module sasic_top (
    input clk,
    input rst_n,
    input in_0,
    input in_1,
    input in_2,
    input in_3,
    input in_4,
    input in_5,
    input in_6,
    input in_7,
    input in_8,
    input in_9,
    input in_10,
    input in_11,
    input in_12,
    input in_13,
    input in_14,
    input in_15,
    input in_16,
    input in_17,
    input in_18,
    input in_19,
    input in_20,
    input in_21,
    input in_22,
    input in_23,
    input in_24,
    input in_25,
    input in_26,
    input in_27,
    input in_28,
    input in_29,
    input in_30,
    input in_31,
    input in_32,
    input in_33,
    input in_34,
    input in_35,
    input in_36,
    input in_37,
    input in_38,
    input in_39,
    output oeb_0,
    output oeb_1,
    output oeb_2,
    output oeb_3,
    output oeb_4,
    output oeb_5,
    output oeb_6,
    output oeb_7,
    output oeb_8,
    output oeb_9,
    output oeb_10,
    output oeb_11,
    output oeb_12,
    output oeb_13,
    output oeb_14,
    output oeb_15,
    output oeb_16,
    output oeb_17,
    output oeb_18,
    output oeb_19,
    output oeb_20,
    output oeb_21,
    output oeb_22,
    output oeb_23,
    output oeb_24,
    output oeb_25,
    output oeb_26,
    output oeb_27,
    output oeb_28,
    output oeb_29,
    output oeb_30,
    output oeb_31,
    output oeb_32,
    output oeb_33,
    output oeb_34,
    output oeb_35,
    output oeb_36,
    output oeb_37,
    output oeb_38,
    output oeb_39,
    output out_0,
    output out_1,
    output out_2,
    output out_3,
    output out_4,
    output out_5,
    output out_6,
    output out_7,
    output out_8,
    output out_9,
    output out_10,
    output out_11,
    output out_12,
    output out_13,
    output out_14,
    output out_15,
    output out_16,
    output out_17,
    output out_18,
    output out_19,
    output out_20,
    output out_21,
    output out_22,
    output out_23,
    output out_24,
    output out_25,
    output out_26,
    output out_27,
    output out_28,
    output out_29,
    output out_30,
    output out_31,
    output out_32,
    output out_33,
    output out_34,
    output out_35,
    output out_36,
    output out_37,
    output out_38,
    output out_39
);

    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9110;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9120;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9132;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9134;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9136;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9138;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9140;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9142;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9160;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9174;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9180;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9182;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9184;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9210;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9226;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9228;
    wire $abc$9276$auto$dfflibmap.cc:532:dfflibmap$9264;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8819;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8821;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8823;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8825;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8827;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8829;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8831;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8833;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8835;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8837;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8839;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8841;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8843;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8845;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8847;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8849;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8851;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8853;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8855;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8857;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8859;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8861;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8863;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8865;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8867;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8869;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8871;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8873;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8875;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8877;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8879;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8881;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8883;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8887;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8889;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8891;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8893;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8895;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8897;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8899;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8901;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8903;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8905;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8907;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8909;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8911;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8913;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8915;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8917;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8921;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8923;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8925;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8927;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8929;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8931;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8933;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8935;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8937;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8939;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8941;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8943;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8945;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8947;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8949;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8951;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8953;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8955;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8957;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8959;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8961;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8963;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8965;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8969;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8971;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8973;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8975;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8979;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8981;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8983;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8987;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8989;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8991;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8993;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8995;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8997;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$8999;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9001;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9003;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9005;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9007;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9009;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9011;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9013;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9015;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9017;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9019;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9021;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9023;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9025;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9027;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9029;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9031;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9033;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9035;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9037;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9039;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9041;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9043;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9045;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9047;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9049;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9051;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9053;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9057;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9061;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9065;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9069;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9073;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9077;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9081;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9085;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9087;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9089;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9091;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9093;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9095;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9097;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9099;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9101;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9103;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9105;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9107;
    wire $abc$9276$auto$rtlil.cc:3205:MuxGate$9109;
    wire $abc$9276$flatten\CPU.$0\adj_bcd[0:0];
    wire $abc$9276$new_n1000;
    wire $abc$9276$new_n1001;
    wire $abc$9276$new_n1002;
    wire $abc$9276$new_n1003;
    wire $abc$9276$new_n1004;
    wire $abc$9276$new_n1005;
    wire $abc$9276$new_n1006;
    wire $abc$9276$new_n1007;
    wire $abc$9276$new_n1008;
    wire $abc$9276$new_n1009;
    wire $abc$9276$new_n1010;
    wire $abc$9276$new_n1011;
    wire $abc$9276$new_n1012;
    wire $abc$9276$new_n1013;
    wire $abc$9276$new_n1014;
    wire $abc$9276$new_n1015;
    wire $abc$9276$new_n1016;
    wire $abc$9276$new_n1017;
    wire $abc$9276$new_n1018;
    wire $abc$9276$new_n1019;
    wire $abc$9276$new_n1020;
    wire $abc$9276$new_n1021;
    wire $abc$9276$new_n1022;
    wire $abc$9276$new_n1023;
    wire $abc$9276$new_n1024;
    wire $abc$9276$new_n1025;
    wire $abc$9276$new_n1026;
    wire $abc$9276$new_n1027;
    wire $abc$9276$new_n1028;
    wire $abc$9276$new_n1029;
    wire $abc$9276$new_n1030;
    wire $abc$9276$new_n1031;
    wire $abc$9276$new_n1032;
    wire $abc$9276$new_n1033;
    wire $abc$9276$new_n1034;
    wire $abc$9276$new_n1035;
    wire $abc$9276$new_n1036;
    wire $abc$9276$new_n1037;
    wire $abc$9276$new_n1039;
    wire $abc$9276$new_n1040;
    wire $abc$9276$new_n1041;
    wire $abc$9276$new_n1042;
    wire $abc$9276$new_n1043;
    wire $abc$9276$new_n1044;
    wire $abc$9276$new_n1045;
    wire $abc$9276$new_n1046;
    wire $abc$9276$new_n1047;
    wire $abc$9276$new_n1048;
    wire $abc$9276$new_n1049;
    wire $abc$9276$new_n1050;
    wire $abc$9276$new_n1051;
    wire $abc$9276$new_n1052;
    wire $abc$9276$new_n1053;
    wire $abc$9276$new_n1054;
    wire $abc$9276$new_n1055;
    wire $abc$9276$new_n1056;
    wire $abc$9276$new_n1058;
    wire $abc$9276$new_n1059;
    wire $abc$9276$new_n1060;
    wire $abc$9276$new_n1061;
    wire $abc$9276$new_n1062;
    wire $abc$9276$new_n1063;
    wire $abc$9276$new_n1064;
    wire $abc$9276$new_n1065;
    wire $abc$9276$new_n1066;
    wire $abc$9276$new_n1067;
    wire $abc$9276$new_n1068;
    wire $abc$9276$new_n1069;
    wire $abc$9276$new_n1070;
    wire $abc$9276$new_n1071;
    wire $abc$9276$new_n1072;
    wire $abc$9276$new_n1073;
    wire $abc$9276$new_n1074;
    wire $abc$9276$new_n1075;
    wire $abc$9276$new_n1076;
    wire $abc$9276$new_n1077;
    wire $abc$9276$new_n1078;
    wire $abc$9276$new_n1079;
    wire $abc$9276$new_n1081;
    wire $abc$9276$new_n1082;
    wire $abc$9276$new_n1083;
    wire $abc$9276$new_n1084;
    wire $abc$9276$new_n1085;
    wire $abc$9276$new_n1086;
    wire $abc$9276$new_n1087;
    wire $abc$9276$new_n1088;
    wire $abc$9276$new_n1089;
    wire $abc$9276$new_n1090;
    wire $abc$9276$new_n1091;
    wire $abc$9276$new_n1092;
    wire $abc$9276$new_n1093;
    wire $abc$9276$new_n1094;
    wire $abc$9276$new_n1095;
    wire $abc$9276$new_n1096;
    wire $abc$9276$new_n1098;
    wire $abc$9276$new_n1099;
    wire $abc$9276$new_n1100;
    wire $abc$9276$new_n1101;
    wire $abc$9276$new_n1102;
    wire $abc$9276$new_n1103;
    wire $abc$9276$new_n1104;
    wire $abc$9276$new_n1105;
    wire $abc$9276$new_n1106;
    wire $abc$9276$new_n1107;
    wire $abc$9276$new_n1108;
    wire $abc$9276$new_n1109;
    wire $abc$9276$new_n1110;
    wire $abc$9276$new_n1111;
    wire $abc$9276$new_n1112;
    wire $abc$9276$new_n1113;
    wire $abc$9276$new_n1115;
    wire $abc$9276$new_n1116;
    wire $abc$9276$new_n1117;
    wire $abc$9276$new_n1118;
    wire $abc$9276$new_n1119;
    wire $abc$9276$new_n1120;
    wire $abc$9276$new_n1121;
    wire $abc$9276$new_n1122;
    wire $abc$9276$new_n1123;
    wire $abc$9276$new_n1124;
    wire $abc$9276$new_n1125;
    wire $abc$9276$new_n1126;
    wire $abc$9276$new_n1127;
    wire $abc$9276$new_n1128;
    wire $abc$9276$new_n1129;
    wire $abc$9276$new_n1130;
    wire $abc$9276$new_n1131;
    wire $abc$9276$new_n1133;
    wire $abc$9276$new_n1134;
    wire $abc$9276$new_n1135;
    wire $abc$9276$new_n1136;
    wire $abc$9276$new_n1137;
    wire $abc$9276$new_n1138;
    wire $abc$9276$new_n1139;
    wire $abc$9276$new_n1140;
    wire $abc$9276$new_n1141;
    wire $abc$9276$new_n1142;
    wire $abc$9276$new_n1143;
    wire $abc$9276$new_n1144;
    wire $abc$9276$new_n1145;
    wire $abc$9276$new_n1146;
    wire $abc$9276$new_n1147;
    wire $abc$9276$new_n1148;
    wire $abc$9276$new_n1150;
    wire $abc$9276$new_n1151;
    wire $abc$9276$new_n1152;
    wire $abc$9276$new_n1153;
    wire $abc$9276$new_n1154;
    wire $abc$9276$new_n1155;
    wire $abc$9276$new_n1156;
    wire $abc$9276$new_n1157;
    wire $abc$9276$new_n1158;
    wire $abc$9276$new_n1159;
    wire $abc$9276$new_n1160;
    wire $abc$9276$new_n1161;
    wire $abc$9276$new_n1162;
    wire $abc$9276$new_n1163;
    wire $abc$9276$new_n1164;
    wire $abc$9276$new_n1165;
    wire $abc$9276$new_n1167;
    wire $abc$9276$new_n1168;
    wire $abc$9276$new_n1169;
    wire $abc$9276$new_n1170;
    wire $abc$9276$new_n1171;
    wire $abc$9276$new_n1172;
    wire $abc$9276$new_n1173;
    wire $abc$9276$new_n1174;
    wire $abc$9276$new_n1175;
    wire $abc$9276$new_n1176;
    wire $abc$9276$new_n1177;
    wire $abc$9276$new_n1178;
    wire $abc$9276$new_n1179;
    wire $abc$9276$new_n1180;
    wire $abc$9276$new_n1181;
    wire $abc$9276$new_n1182;
    wire $abc$9276$new_n1183;
    wire $abc$9276$new_n1184;
    wire $abc$9276$new_n1185;
    wire $abc$9276$new_n1187;
    wire $abc$9276$new_n1188;
    wire $abc$9276$new_n1189;
    wire $abc$9276$new_n1190;
    wire $abc$9276$new_n1191;
    wire $abc$9276$new_n1192;
    wire $abc$9276$new_n1193;
    wire $abc$9276$new_n1194;
    wire $abc$9276$new_n1195;
    wire $abc$9276$new_n1196;
    wire $abc$9276$new_n1197;
    wire $abc$9276$new_n1198;
    wire $abc$9276$new_n1199;
    wire $abc$9276$new_n1200;
    wire $abc$9276$new_n1201;
    wire $abc$9276$new_n1202;
    wire $abc$9276$new_n1203;
    wire $abc$9276$new_n1204;
    wire $abc$9276$new_n1206;
    wire $abc$9276$new_n1207;
    wire $abc$9276$new_n1208;
    wire $abc$9276$new_n1209;
    wire $abc$9276$new_n1210;
    wire $abc$9276$new_n1211;
    wire $abc$9276$new_n1212;
    wire $abc$9276$new_n1213;
    wire $abc$9276$new_n1214;
    wire $abc$9276$new_n1215;
    wire $abc$9276$new_n1216;
    wire $abc$9276$new_n1217;
    wire $abc$9276$new_n1218;
    wire $abc$9276$new_n1219;
    wire $abc$9276$new_n1220;
    wire $abc$9276$new_n1221;
    wire $abc$9276$new_n1222;
    wire $abc$9276$new_n1223;
    wire $abc$9276$new_n1224;
    wire $abc$9276$new_n1226;
    wire $abc$9276$new_n1227;
    wire $abc$9276$new_n1228;
    wire $abc$9276$new_n1229;
    wire $abc$9276$new_n1230;
    wire $abc$9276$new_n1231;
    wire $abc$9276$new_n1232;
    wire $abc$9276$new_n1233;
    wire $abc$9276$new_n1234;
    wire $abc$9276$new_n1235;
    wire $abc$9276$new_n1236;
    wire $abc$9276$new_n1237;
    wire $abc$9276$new_n1238;
    wire $abc$9276$new_n1239;
    wire $abc$9276$new_n1240;
    wire $abc$9276$new_n1241;
    wire $abc$9276$new_n1242;
    wire $abc$9276$new_n1243;
    wire $abc$9276$new_n1245;
    wire $abc$9276$new_n1246;
    wire $abc$9276$new_n1247;
    wire $abc$9276$new_n1248;
    wire $abc$9276$new_n1249;
    wire $abc$9276$new_n1250;
    wire $abc$9276$new_n1251;
    wire $abc$9276$new_n1252;
    wire $abc$9276$new_n1253;
    wire $abc$9276$new_n1254;
    wire $abc$9276$new_n1255;
    wire $abc$9276$new_n1256;
    wire $abc$9276$new_n1257;
    wire $abc$9276$new_n1258;
    wire $abc$9276$new_n1259;
    wire $abc$9276$new_n1260;
    wire $abc$9276$new_n1261;
    wire $abc$9276$new_n1262;
    wire $abc$9276$new_n1263;
    wire $abc$9276$new_n1264;
    wire $abc$9276$new_n1266;
    wire $abc$9276$new_n1267;
    wire $abc$9276$new_n1268;
    wire $abc$9276$new_n1269;
    wire $abc$9276$new_n1270;
    wire $abc$9276$new_n1271;
    wire $abc$9276$new_n1272;
    wire $abc$9276$new_n1273;
    wire $abc$9276$new_n1274;
    wire $abc$9276$new_n1275;
    wire $abc$9276$new_n1276;
    wire $abc$9276$new_n1277;
    wire $abc$9276$new_n1278;
    wire $abc$9276$new_n1279;
    wire $abc$9276$new_n1280;
    wire $abc$9276$new_n1281;
    wire $abc$9276$new_n1282;
    wire $abc$9276$new_n1283;
    wire $abc$9276$new_n1284;
    wire $abc$9276$new_n1286;
    wire $abc$9276$new_n1287;
    wire $abc$9276$new_n1288;
    wire $abc$9276$new_n1289;
    wire $abc$9276$new_n1290;
    wire $abc$9276$new_n1291;
    wire $abc$9276$new_n1292;
    wire $abc$9276$new_n1293;
    wire $abc$9276$new_n1294;
    wire $abc$9276$new_n1295;
    wire $abc$9276$new_n1296;
    wire $abc$9276$new_n1297;
    wire $abc$9276$new_n1298;
    wire $abc$9276$new_n1299;
    wire $abc$9276$new_n1300;
    wire $abc$9276$new_n1301;
    wire $abc$9276$new_n1302;
    wire $abc$9276$new_n1304;
    wire $abc$9276$new_n1305;
    wire $abc$9276$new_n1306;
    wire $abc$9276$new_n1307;
    wire $abc$9276$new_n1308;
    wire $abc$9276$new_n1309;
    wire $abc$9276$new_n1310;
    wire $abc$9276$new_n1311;
    wire $abc$9276$new_n1312;
    wire $abc$9276$new_n1313;
    wire $abc$9276$new_n1314;
    wire $abc$9276$new_n1315;
    wire $abc$9276$new_n1316;
    wire $abc$9276$new_n1317;
    wire $abc$9276$new_n1318;
    wire $abc$9276$new_n1319;
    wire $abc$9276$new_n1321;
    wire $abc$9276$new_n1322;
    wire $abc$9276$new_n1324;
    wire $abc$9276$new_n1325;
    wire $abc$9276$new_n1327;
    wire $abc$9276$new_n1328;
    wire $abc$9276$new_n1330;
    wire $abc$9276$new_n1331;
    wire $abc$9276$new_n1332;
    wire $abc$9276$new_n1333;
    wire $abc$9276$new_n1334;
    wire $abc$9276$new_n1335;
    wire $abc$9276$new_n1336;
    wire $abc$9276$new_n1337;
    wire $abc$9276$new_n1338;
    wire $abc$9276$new_n1339;
    wire $abc$9276$new_n1340;
    wire $abc$9276$new_n1341;
    wire $abc$9276$new_n1342;
    wire $abc$9276$new_n1343;
    wire $abc$9276$new_n1344;
    wire $abc$9276$new_n1345;
    wire $abc$9276$new_n1347;
    wire $abc$9276$new_n1348;
    wire $abc$9276$new_n1349;
    wire $abc$9276$new_n1350;
    wire $abc$9276$new_n1351;
    wire $abc$9276$new_n1352;
    wire $abc$9276$new_n1353;
    wire $abc$9276$new_n1354;
    wire $abc$9276$new_n1355;
    wire $abc$9276$new_n1356;
    wire $abc$9276$new_n1357;
    wire $abc$9276$new_n1358;
    wire $abc$9276$new_n1359;
    wire $abc$9276$new_n1360;
    wire $abc$9276$new_n1361;
    wire $abc$9276$new_n1362;
    wire $abc$9276$new_n1363;
    wire $abc$9276$new_n1364;
    wire $abc$9276$new_n1366;
    wire $abc$9276$new_n1367;
    wire $abc$9276$new_n1368;
    wire $abc$9276$new_n1369;
    wire $abc$9276$new_n1370;
    wire $abc$9276$new_n1371;
    wire $abc$9276$new_n1372;
    wire $abc$9276$new_n1373;
    wire $abc$9276$new_n1374;
    wire $abc$9276$new_n1375;
    wire $abc$9276$new_n1376;
    wire $abc$9276$new_n1377;
    wire $abc$9276$new_n1378;
    wire $abc$9276$new_n1379;
    wire $abc$9276$new_n1380;
    wire $abc$9276$new_n1381;
    wire $abc$9276$new_n1382;
    wire $abc$9276$new_n1383;
    wire $abc$9276$new_n1384;
    wire $abc$9276$new_n1385;
    wire $abc$9276$new_n1386;
    wire $abc$9276$new_n1387;
    wire $abc$9276$new_n1388;
    wire $abc$9276$new_n1389;
    wire $abc$9276$new_n1390;
    wire $abc$9276$new_n1392;
    wire $abc$9276$new_n1393;
    wire $abc$9276$new_n1394;
    wire $abc$9276$new_n1395;
    wire $abc$9276$new_n1396;
    wire $abc$9276$new_n1397;
    wire $abc$9276$new_n1398;
    wire $abc$9276$new_n1399;
    wire $abc$9276$new_n1400;
    wire $abc$9276$new_n1401;
    wire $abc$9276$new_n1402;
    wire $abc$9276$new_n1403;
    wire $abc$9276$new_n1404;
    wire $abc$9276$new_n1405;
    wire $abc$9276$new_n1406;
    wire $abc$9276$new_n1407;
    wire $abc$9276$new_n1408;
    wire $abc$9276$new_n1409;
    wire $abc$9276$new_n1410;
    wire $abc$9276$new_n1411;
    wire $abc$9276$new_n1412;
    wire $abc$9276$new_n1413;
    wire $abc$9276$new_n1414;
    wire $abc$9276$new_n1415;
    wire $abc$9276$new_n1416;
    wire $abc$9276$new_n1417;
    wire $abc$9276$new_n1418;
    wire $abc$9276$new_n1419;
    wire $abc$9276$new_n1420;
    wire $abc$9276$new_n1421;
    wire $abc$9276$new_n1422;
    wire $abc$9276$new_n1423;
    wire $abc$9276$new_n1424;
    wire $abc$9276$new_n1426;
    wire $abc$9276$new_n1428;
    wire $abc$9276$new_n1429;
    wire $abc$9276$new_n1430;
    wire $abc$9276$new_n1431;
    wire $abc$9276$new_n1432;
    wire $abc$9276$new_n1433;
    wire $abc$9276$new_n1434;
    wire $abc$9276$new_n1435;
    wire $abc$9276$new_n1436;
    wire $abc$9276$new_n1437;
    wire $abc$9276$new_n1438;
    wire $abc$9276$new_n1439;
    wire $abc$9276$new_n1440;
    wire $abc$9276$new_n1441;
    wire $abc$9276$new_n1442;
    wire $abc$9276$new_n1443;
    wire $abc$9276$new_n1444;
    wire $abc$9276$new_n1445;
    wire $abc$9276$new_n1446;
    wire $abc$9276$new_n1447;
    wire $abc$9276$new_n1448;
    wire $abc$9276$new_n1449;
    wire $abc$9276$new_n1450;
    wire $abc$9276$new_n1451;
    wire $abc$9276$new_n1452;
    wire $abc$9276$new_n1453;
    wire $abc$9276$new_n1454;
    wire $abc$9276$new_n1455;
    wire $abc$9276$new_n1456;
    wire $abc$9276$new_n1457;
    wire $abc$9276$new_n1458;
    wire $abc$9276$new_n1459;
    wire $abc$9276$new_n1460;
    wire $abc$9276$new_n1461;
    wire $abc$9276$new_n1462;
    wire $abc$9276$new_n1463;
    wire $abc$9276$new_n1464;
    wire $abc$9276$new_n1465;
    wire $abc$9276$new_n1466;
    wire $abc$9276$new_n1467;
    wire $abc$9276$new_n1468;
    wire $abc$9276$new_n1469;
    wire $abc$9276$new_n1470;
    wire $abc$9276$new_n1471;
    wire $abc$9276$new_n1472;
    wire $abc$9276$new_n1473;
    wire $abc$9276$new_n1474;
    wire $abc$9276$new_n1475;
    wire $abc$9276$new_n1476;
    wire $abc$9276$new_n1477;
    wire $abc$9276$new_n1478;
    wire $abc$9276$new_n1479;
    wire $abc$9276$new_n1480;
    wire $abc$9276$new_n1481;
    wire $abc$9276$new_n1482;
    wire $abc$9276$new_n1483;
    wire $abc$9276$new_n1484;
    wire $abc$9276$new_n1485;
    wire $abc$9276$new_n1486;
    wire $abc$9276$new_n1487;
    wire $abc$9276$new_n1488;
    wire $abc$9276$new_n1489;
    wire $abc$9276$new_n1490;
    wire $abc$9276$new_n1491;
    wire $abc$9276$new_n1492;
    wire $abc$9276$new_n1493;
    wire $abc$9276$new_n1494;
    wire $abc$9276$new_n1495;
    wire $abc$9276$new_n1496;
    wire $abc$9276$new_n1497;
    wire $abc$9276$new_n1498;
    wire $abc$9276$new_n1499;
    wire $abc$9276$new_n1500;
    wire $abc$9276$new_n1502;
    wire $abc$9276$new_n1503;
    wire $abc$9276$new_n1504;
    wire $abc$9276$new_n1505;
    wire $abc$9276$new_n1506;
    wire $abc$9276$new_n1507;
    wire $abc$9276$new_n1508;
    wire $abc$9276$new_n1509;
    wire $abc$9276$new_n1510;
    wire $abc$9276$new_n1511;
    wire $abc$9276$new_n1513;
    wire $abc$9276$new_n1514;
    wire $abc$9276$new_n1515;
    wire $abc$9276$new_n1516;
    wire $abc$9276$new_n1517;
    wire $abc$9276$new_n1518;
    wire $abc$9276$new_n1519;
    wire $abc$9276$new_n1520;
    wire $abc$9276$new_n1521;
    wire $abc$9276$new_n1522;
    wire $abc$9276$new_n1523;
    wire $abc$9276$new_n1524;
    wire $abc$9276$new_n1525;
    wire $abc$9276$new_n1526;
    wire $abc$9276$new_n1527;
    wire $abc$9276$new_n1528;
    wire $abc$9276$new_n1529;
    wire $abc$9276$new_n1530;
    wire $abc$9276$new_n1531;
    wire $abc$9276$new_n1533;
    wire $abc$9276$new_n1534;
    wire $abc$9276$new_n1536;
    wire $abc$9276$new_n1537;
    wire $abc$9276$new_n1538;
    wire $abc$9276$new_n1539;
    wire $abc$9276$new_n1540;
    wire $abc$9276$new_n1541;
    wire $abc$9276$new_n1542;
    wire $abc$9276$new_n1543;
    wire $abc$9276$new_n1544;
    wire $abc$9276$new_n1545;
    wire $abc$9276$new_n1546;
    wire $abc$9276$new_n1547;
    wire $abc$9276$new_n1548;
    wire $abc$9276$new_n1549;
    wire $abc$9276$new_n1550;
    wire $abc$9276$new_n1551;
    wire $abc$9276$new_n1552;
    wire $abc$9276$new_n1553;
    wire $abc$9276$new_n1554;
    wire $abc$9276$new_n1555;
    wire $abc$9276$new_n1556;
    wire $abc$9276$new_n1558;
    wire $abc$9276$new_n1559;
    wire $abc$9276$new_n1561;
    wire $abc$9276$new_n1562;
    wire $abc$9276$new_n1563;
    wire $abc$9276$new_n1564;
    wire $abc$9276$new_n1565;
    wire $abc$9276$new_n1566;
    wire $abc$9276$new_n1567;
    wire $abc$9276$new_n1568;
    wire $abc$9276$new_n1569;
    wire $abc$9276$new_n1570;
    wire $abc$9276$new_n1571;
    wire $abc$9276$new_n1572;
    wire $abc$9276$new_n1573;
    wire $abc$9276$new_n1574;
    wire $abc$9276$new_n1575;
    wire $abc$9276$new_n1576;
    wire $abc$9276$new_n1577;
    wire $abc$9276$new_n1578;
    wire $abc$9276$new_n1579;
    wire $abc$9276$new_n1580;
    wire $abc$9276$new_n1581;
    wire $abc$9276$new_n1582;
    wire $abc$9276$new_n1584;
    wire $abc$9276$new_n1585;
    wire $abc$9276$new_n1587;
    wire $abc$9276$new_n1588;
    wire $abc$9276$new_n1589;
    wire $abc$9276$new_n1590;
    wire $abc$9276$new_n1591;
    wire $abc$9276$new_n1592;
    wire $abc$9276$new_n1593;
    wire $abc$9276$new_n1594;
    wire $abc$9276$new_n1595;
    wire $abc$9276$new_n1596;
    wire $abc$9276$new_n1597;
    wire $abc$9276$new_n1598;
    wire $abc$9276$new_n1599;
    wire $abc$9276$new_n1600;
    wire $abc$9276$new_n1601;
    wire $abc$9276$new_n1602;
    wire $abc$9276$new_n1603;
    wire $abc$9276$new_n1604;
    wire $abc$9276$new_n1605;
    wire $abc$9276$new_n1606;
    wire $abc$9276$new_n1607;
    wire $abc$9276$new_n1608;
    wire $abc$9276$new_n1610;
    wire $abc$9276$new_n1611;
    wire $abc$9276$new_n1613;
    wire $abc$9276$new_n1614;
    wire $abc$9276$new_n1615;
    wire $abc$9276$new_n1616;
    wire $abc$9276$new_n1617;
    wire $abc$9276$new_n1618;
    wire $abc$9276$new_n1619;
    wire $abc$9276$new_n1620;
    wire $abc$9276$new_n1621;
    wire $abc$9276$new_n1622;
    wire $abc$9276$new_n1623;
    wire $abc$9276$new_n1624;
    wire $abc$9276$new_n1625;
    wire $abc$9276$new_n1626;
    wire $abc$9276$new_n1627;
    wire $abc$9276$new_n1628;
    wire $abc$9276$new_n1629;
    wire $abc$9276$new_n1630;
    wire $abc$9276$new_n1631;
    wire $abc$9276$new_n1632;
    wire $abc$9276$new_n1633;
    wire $abc$9276$new_n1634;
    wire $abc$9276$new_n1636;
    wire $abc$9276$new_n1637;
    wire $abc$9276$new_n1639;
    wire $abc$9276$new_n1640;
    wire $abc$9276$new_n1641;
    wire $abc$9276$new_n1642;
    wire $abc$9276$new_n1643;
    wire $abc$9276$new_n1644;
    wire $abc$9276$new_n1645;
    wire $abc$9276$new_n1646;
    wire $abc$9276$new_n1647;
    wire $abc$9276$new_n1648;
    wire $abc$9276$new_n1649;
    wire $abc$9276$new_n1650;
    wire $abc$9276$new_n1651;
    wire $abc$9276$new_n1652;
    wire $abc$9276$new_n1653;
    wire $abc$9276$new_n1654;
    wire $abc$9276$new_n1655;
    wire $abc$9276$new_n1656;
    wire $abc$9276$new_n1657;
    wire $abc$9276$new_n1658;
    wire $abc$9276$new_n1659;
    wire $abc$9276$new_n1660;
    wire $abc$9276$new_n1662;
    wire $abc$9276$new_n1663;
    wire $abc$9276$new_n1665;
    wire $abc$9276$new_n1666;
    wire $abc$9276$new_n1667;
    wire $abc$9276$new_n1668;
    wire $abc$9276$new_n1669;
    wire $abc$9276$new_n1670;
    wire $abc$9276$new_n1671;
    wire $abc$9276$new_n1672;
    wire $abc$9276$new_n1673;
    wire $abc$9276$new_n1674;
    wire $abc$9276$new_n1675;
    wire $abc$9276$new_n1676;
    wire $abc$9276$new_n1677;
    wire $abc$9276$new_n1678;
    wire $abc$9276$new_n1679;
    wire $abc$9276$new_n1680;
    wire $abc$9276$new_n1681;
    wire $abc$9276$new_n1682;
    wire $abc$9276$new_n1683;
    wire $abc$9276$new_n1684;
    wire $abc$9276$new_n1686;
    wire $abc$9276$new_n1687;
    wire $abc$9276$new_n1689;
    wire $abc$9276$new_n1690;
    wire $abc$9276$new_n1691;
    wire $abc$9276$new_n1692;
    wire $abc$9276$new_n1693;
    wire $abc$9276$new_n1694;
    wire $abc$9276$new_n1695;
    wire $abc$9276$new_n1696;
    wire $abc$9276$new_n1697;
    wire $abc$9276$new_n1698;
    wire $abc$9276$new_n1700;
    wire $abc$9276$new_n1701;
    wire $abc$9276$new_n1703;
    wire $abc$9276$new_n1704;
    wire $abc$9276$new_n1705;
    wire $abc$9276$new_n1706;
    wire $abc$9276$new_n1707;
    wire $abc$9276$new_n1708;
    wire $abc$9276$new_n1709;
    wire $abc$9276$new_n1710;
    wire $abc$9276$new_n1712;
    wire $abc$9276$new_n1713;
    wire $abc$9276$new_n1715;
    wire $abc$9276$new_n1716;
    wire $abc$9276$new_n1717;
    wire $abc$9276$new_n1718;
    wire $abc$9276$new_n1719;
    wire $abc$9276$new_n1720;
    wire $abc$9276$new_n1721;
    wire $abc$9276$new_n1722;
    wire $abc$9276$new_n1724;
    wire $abc$9276$new_n1725;
    wire $abc$9276$new_n1727;
    wire $abc$9276$new_n1728;
    wire $abc$9276$new_n1729;
    wire $abc$9276$new_n1730;
    wire $abc$9276$new_n1731;
    wire $abc$9276$new_n1732;
    wire $abc$9276$new_n1733;
    wire $abc$9276$new_n1734;
    wire $abc$9276$new_n1736;
    wire $abc$9276$new_n1737;
    wire $abc$9276$new_n1739;
    wire $abc$9276$new_n1740;
    wire $abc$9276$new_n1741;
    wire $abc$9276$new_n1742;
    wire $abc$9276$new_n1743;
    wire $abc$9276$new_n1744;
    wire $abc$9276$new_n1745;
    wire $abc$9276$new_n1746;
    wire $abc$9276$new_n1748;
    wire $abc$9276$new_n1749;
    wire $abc$9276$new_n1751;
    wire $abc$9276$new_n1752;
    wire $abc$9276$new_n1753;
    wire $abc$9276$new_n1754;
    wire $abc$9276$new_n1755;
    wire $abc$9276$new_n1756;
    wire $abc$9276$new_n1757;
    wire $abc$9276$new_n1758;
    wire $abc$9276$new_n1760;
    wire $abc$9276$new_n1761;
    wire $abc$9276$new_n1763;
    wire $abc$9276$new_n1764;
    wire $abc$9276$new_n1765;
    wire $abc$9276$new_n1766;
    wire $abc$9276$new_n1767;
    wire $abc$9276$new_n1768;
    wire $abc$9276$new_n1769;
    wire $abc$9276$new_n1770;
    wire $abc$9276$new_n1771;
    wire $abc$9276$new_n1772;
    wire $abc$9276$new_n1774;
    wire $abc$9276$new_n1775;
    wire $abc$9276$new_n1777;
    wire $abc$9276$new_n1778;
    wire $abc$9276$new_n1779;
    wire $abc$9276$new_n1780;
    wire $abc$9276$new_n1781;
    wire $abc$9276$new_n1782;
    wire $abc$9276$new_n1783;
    wire $abc$9276$new_n1784;
    wire $abc$9276$new_n1786;
    wire $abc$9276$new_n1787;
    wire $abc$9276$new_n1789;
    wire $abc$9276$new_n1790;
    wire $abc$9276$new_n1791;
    wire $abc$9276$new_n1792;
    wire $abc$9276$new_n1793;
    wire $abc$9276$new_n1795;
    wire $abc$9276$new_n1796;
    wire $abc$9276$new_n1798;
    wire $abc$9276$new_n1799;
    wire $abc$9276$new_n1801;
    wire $abc$9276$new_n1802;
    wire $abc$9276$new_n1804;
    wire $abc$9276$new_n1805;
    wire $abc$9276$new_n1807;
    wire $abc$9276$new_n1808;
    wire $abc$9276$new_n1810;
    wire $abc$9276$new_n1811;
    wire $abc$9276$new_n1813;
    wire $abc$9276$new_n1814;
    wire $abc$9276$new_n1816;
    wire $abc$9276$new_n1817;
    wire $abc$9276$new_n1818;
    wire $abc$9276$new_n1819;
    wire $abc$9276$new_n1820;
    wire $abc$9276$new_n1821;
    wire $abc$9276$new_n1822;
    wire $abc$9276$new_n1823;
    wire $abc$9276$new_n1824;
    wire $abc$9276$new_n1825;
    wire $abc$9276$new_n1826;
    wire $abc$9276$new_n1827;
    wire $abc$9276$new_n1828;
    wire $abc$9276$new_n1829;
    wire $abc$9276$new_n1830;
    wire $abc$9276$new_n1831;
    wire $abc$9276$new_n1832;
    wire $abc$9276$new_n1833;
    wire $abc$9276$new_n1834;
    wire $abc$9276$new_n1835;
    wire $abc$9276$new_n1836;
    wire $abc$9276$new_n1837;
    wire $abc$9276$new_n1838;
    wire $abc$9276$new_n1839;
    wire $abc$9276$new_n1840;
    wire $abc$9276$new_n1841;
    wire $abc$9276$new_n1842;
    wire $abc$9276$new_n1843;
    wire $abc$9276$new_n1844;
    wire $abc$9276$new_n1845;
    wire $abc$9276$new_n1846;
    wire $abc$9276$new_n1847;
    wire $abc$9276$new_n1848;
    wire $abc$9276$new_n1849;
    wire $abc$9276$new_n1850;
    wire $abc$9276$new_n1851;
    wire $abc$9276$new_n1852;
    wire $abc$9276$new_n1853;
    wire $abc$9276$new_n1854;
    wire $abc$9276$new_n1855;
    wire $abc$9276$new_n1856;
    wire $abc$9276$new_n1857;
    wire $abc$9276$new_n1858;
    wire $abc$9276$new_n1859;
    wire $abc$9276$new_n1860;
    wire $abc$9276$new_n1861;
    wire $abc$9276$new_n1862;
    wire $abc$9276$new_n1863;
    wire $abc$9276$new_n1864;
    wire $abc$9276$new_n1865;
    wire $abc$9276$new_n1866;
    wire $abc$9276$new_n1867;
    wire $abc$9276$new_n1868;
    wire $abc$9276$new_n1869;
    wire $abc$9276$new_n1870;
    wire $abc$9276$new_n1871;
    wire $abc$9276$new_n1872;
    wire $abc$9276$new_n1873;
    wire $abc$9276$new_n1874;
    wire $abc$9276$new_n1875;
    wire $abc$9276$new_n1876;
    wire $abc$9276$new_n1877;
    wire $abc$9276$new_n1878;
    wire $abc$9276$new_n1879;
    wire $abc$9276$new_n1880;
    wire $abc$9276$new_n1881;
    wire $abc$9276$new_n1882;
    wire $abc$9276$new_n1883;
    wire $abc$9276$new_n1884;
    wire $abc$9276$new_n1885;
    wire $abc$9276$new_n1886;
    wire $abc$9276$new_n1887;
    wire $abc$9276$new_n1888;
    wire $abc$9276$new_n1889;
    wire $abc$9276$new_n1890;
    wire $abc$9276$new_n1891;
    wire $abc$9276$new_n1892;
    wire $abc$9276$new_n1893;
    wire $abc$9276$new_n1894;
    wire $abc$9276$new_n1895;
    wire $abc$9276$new_n1896;
    wire $abc$9276$new_n1897;
    wire $abc$9276$new_n1898;
    wire $abc$9276$new_n1899;
    wire $abc$9276$new_n1900;
    wire $abc$9276$new_n1901;
    wire $abc$9276$new_n1902;
    wire $abc$9276$new_n1903;
    wire $abc$9276$new_n1904;
    wire $abc$9276$new_n1905;
    wire $abc$9276$new_n1906;
    wire $abc$9276$new_n1907;
    wire $abc$9276$new_n1908;
    wire $abc$9276$new_n1909;
    wire $abc$9276$new_n1910;
    wire $abc$9276$new_n1911;
    wire $abc$9276$new_n1912;
    wire $abc$9276$new_n1913;
    wire $abc$9276$new_n1914;
    wire $abc$9276$new_n1915;
    wire $abc$9276$new_n1916;
    wire $abc$9276$new_n1917;
    wire $abc$9276$new_n1918;
    wire $abc$9276$new_n1919;
    wire $abc$9276$new_n1920;
    wire $abc$9276$new_n1921;
    wire $abc$9276$new_n1922;
    wire $abc$9276$new_n1923;
    wire $abc$9276$new_n1924;
    wire $abc$9276$new_n1925;
    wire $abc$9276$new_n1926;
    wire $abc$9276$new_n1927;
    wire $abc$9276$new_n1928;
    wire $abc$9276$new_n1929;
    wire $abc$9276$new_n1930;
    wire $abc$9276$new_n1931;
    wire $abc$9276$new_n1932;
    wire $abc$9276$new_n1933;
    wire $abc$9276$new_n1934;
    wire $abc$9276$new_n1935;
    wire $abc$9276$new_n1936;
    wire $abc$9276$new_n1937;
    wire $abc$9276$new_n1938;
    wire $abc$9276$new_n1939;
    wire $abc$9276$new_n1940;
    wire $abc$9276$new_n1941;
    wire $abc$9276$new_n1942;
    wire $abc$9276$new_n1943;
    wire $abc$9276$new_n1945;
    wire $abc$9276$new_n1946;
    wire $abc$9276$new_n1947;
    wire $abc$9276$new_n1948;
    wire $abc$9276$new_n1949;
    wire $abc$9276$new_n1950;
    wire $abc$9276$new_n1951;
    wire $abc$9276$new_n1952;
    wire $abc$9276$new_n1953;
    wire $abc$9276$new_n1954;
    wire $abc$9276$new_n1955;
    wire $abc$9276$new_n1956;
    wire $abc$9276$new_n1957;
    wire $abc$9276$new_n1958;
    wire $abc$9276$new_n1959;
    wire $abc$9276$new_n1960;
    wire $abc$9276$new_n1961;
    wire $abc$9276$new_n1962;
    wire $abc$9276$new_n1963;
    wire $abc$9276$new_n1964;
    wire $abc$9276$new_n1965;
    wire $abc$9276$new_n1966;
    wire $abc$9276$new_n1967;
    wire $abc$9276$new_n1968;
    wire $abc$9276$new_n1969;
    wire $abc$9276$new_n1970;
    wire $abc$9276$new_n1971;
    wire $abc$9276$new_n1972;
    wire $abc$9276$new_n1973;
    wire $abc$9276$new_n1974;
    wire $abc$9276$new_n1975;
    wire $abc$9276$new_n1976;
    wire $abc$9276$new_n1977;
    wire $abc$9276$new_n1978;
    wire $abc$9276$new_n1979;
    wire $abc$9276$new_n1980;
    wire $abc$9276$new_n1981;
    wire $abc$9276$new_n1982;
    wire $abc$9276$new_n1983;
    wire $abc$9276$new_n1984;
    wire $abc$9276$new_n1985;
    wire $abc$9276$new_n1986;
    wire $abc$9276$new_n1987;
    wire $abc$9276$new_n1988;
    wire $abc$9276$new_n1989;
    wire $abc$9276$new_n1990;
    wire $abc$9276$new_n1991;
    wire $abc$9276$new_n1992;
    wire $abc$9276$new_n1993;
    wire $abc$9276$new_n1994;
    wire $abc$9276$new_n1995;
    wire $abc$9276$new_n1996;
    wire $abc$9276$new_n1997;
    wire $abc$9276$new_n1998;
    wire $abc$9276$new_n2000;
    wire $abc$9276$new_n2001;
    wire $abc$9276$new_n2002;
    wire $abc$9276$new_n2003;
    wire $abc$9276$new_n2004;
    wire $abc$9276$new_n2005;
    wire $abc$9276$new_n2006;
    wire $abc$9276$new_n2007;
    wire $abc$9276$new_n2008;
    wire $abc$9276$new_n2009;
    wire $abc$9276$new_n2010;
    wire $abc$9276$new_n2011;
    wire $abc$9276$new_n2012;
    wire $abc$9276$new_n2013;
    wire $abc$9276$new_n2014;
    wire $abc$9276$new_n2015;
    wire $abc$9276$new_n2016;
    wire $abc$9276$new_n2017;
    wire $abc$9276$new_n2018;
    wire $abc$9276$new_n2019;
    wire $abc$9276$new_n2020;
    wire $abc$9276$new_n2021;
    wire $abc$9276$new_n2022;
    wire $abc$9276$new_n2024;
    wire $abc$9276$new_n2025;
    wire $abc$9276$new_n2026;
    wire $abc$9276$new_n2027;
    wire $abc$9276$new_n2028;
    wire $abc$9276$new_n2029;
    wire $abc$9276$new_n2030;
    wire $abc$9276$new_n2031;
    wire $abc$9276$new_n2032;
    wire $abc$9276$new_n2033;
    wire $abc$9276$new_n2034;
    wire $abc$9276$new_n2035;
    wire $abc$9276$new_n2036;
    wire $abc$9276$new_n2037;
    wire $abc$9276$new_n2038;
    wire $abc$9276$new_n2039;
    wire $abc$9276$new_n2040;
    wire $abc$9276$new_n2041;
    wire $abc$9276$new_n2042;
    wire $abc$9276$new_n2043;
    wire $abc$9276$new_n2044;
    wire $abc$9276$new_n2045;
    wire $abc$9276$new_n2046;
    wire $abc$9276$new_n2047;
    wire $abc$9276$new_n2048;
    wire $abc$9276$new_n2049;
    wire $abc$9276$new_n2051;
    wire $abc$9276$new_n2052;
    wire $abc$9276$new_n2053;
    wire $abc$9276$new_n2054;
    wire $abc$9276$new_n2055;
    wire $abc$9276$new_n2056;
    wire $abc$9276$new_n2057;
    wire $abc$9276$new_n2058;
    wire $abc$9276$new_n2059;
    wire $abc$9276$new_n2060;
    wire $abc$9276$new_n2061;
    wire $abc$9276$new_n2062;
    wire $abc$9276$new_n2063;
    wire $abc$9276$new_n2064;
    wire $abc$9276$new_n2065;
    wire $abc$9276$new_n2066;
    wire $abc$9276$new_n2067;
    wire $abc$9276$new_n2068;
    wire $abc$9276$new_n2070;
    wire $abc$9276$new_n2071;
    wire $abc$9276$new_n2072;
    wire $abc$9276$new_n2073;
    wire $abc$9276$new_n2074;
    wire $abc$9276$new_n2075;
    wire $abc$9276$new_n2076;
    wire $abc$9276$new_n2077;
    wire $abc$9276$new_n2078;
    wire $abc$9276$new_n2079;
    wire $abc$9276$new_n2080;
    wire $abc$9276$new_n2081;
    wire $abc$9276$new_n2082;
    wire $abc$9276$new_n2084;
    wire $abc$9276$new_n2085;
    wire $abc$9276$new_n2086;
    wire $abc$9276$new_n2087;
    wire $abc$9276$new_n2088;
    wire $abc$9276$new_n2089;
    wire $abc$9276$new_n2090;
    wire $abc$9276$new_n2091;
    wire $abc$9276$new_n2092;
    wire $abc$9276$new_n2093;
    wire $abc$9276$new_n2094;
    wire $abc$9276$new_n2095;
    wire $abc$9276$new_n2096;
    wire $abc$9276$new_n2097;
    wire $abc$9276$new_n2098;
    wire $abc$9276$new_n2100;
    wire $abc$9276$new_n2101;
    wire $abc$9276$new_n2102;
    wire $abc$9276$new_n2103;
    wire $abc$9276$new_n2104;
    wire $abc$9276$new_n2105;
    wire $abc$9276$new_n2106;
    wire $abc$9276$new_n2107;
    wire $abc$9276$new_n2109;
    wire $abc$9276$new_n2110;
    wire $abc$9276$new_n2111;
    wire $abc$9276$new_n2112;
    wire $abc$9276$new_n2113;
    wire $abc$9276$new_n2114;
    wire $abc$9276$new_n2115;
    wire $abc$9276$new_n2116;
    wire $abc$9276$new_n2117;
    wire $abc$9276$new_n2118;
    wire $abc$9276$new_n2119;
    wire $abc$9276$new_n2120;
    wire $abc$9276$new_n2121;
    wire $abc$9276$new_n2122;
    wire $abc$9276$new_n2123;
    wire $abc$9276$new_n2124;
    wire $abc$9276$new_n2125;
    wire $abc$9276$new_n2127;
    wire $abc$9276$new_n2128;
    wire $abc$9276$new_n2129;
    wire $abc$9276$new_n2130;
    wire $abc$9276$new_n2131;
    wire $abc$9276$new_n2133;
    wire $abc$9276$new_n2134;
    wire $abc$9276$new_n2135;
    wire $abc$9276$new_n2136;
    wire $abc$9276$new_n2137;
    wire $abc$9276$new_n2138;
    wire $abc$9276$new_n2139;
    wire $abc$9276$new_n2140;
    wire $abc$9276$new_n2141;
    wire $abc$9276$new_n2142;
    wire $abc$9276$new_n2143;
    wire $abc$9276$new_n2144;
    wire $abc$9276$new_n2145;
    wire $abc$9276$new_n2147;
    wire $abc$9276$new_n2148;
    wire $abc$9276$new_n2149;
    wire $abc$9276$new_n2150;
    wire $abc$9276$new_n2151;
    wire $abc$9276$new_n2152;
    wire $abc$9276$new_n2153;
    wire $abc$9276$new_n2154;
    wire $abc$9276$new_n2155;
    wire $abc$9276$new_n2156;
    wire $abc$9276$new_n2157;
    wire $abc$9276$new_n2158;
    wire $abc$9276$new_n2160;
    wire $abc$9276$new_n2161;
    wire $abc$9276$new_n2162;
    wire $abc$9276$new_n2163;
    wire $abc$9276$new_n2164;
    wire $abc$9276$new_n2165;
    wire $abc$9276$new_n2166;
    wire $abc$9276$new_n2167;
    wire $abc$9276$new_n2168;
    wire $abc$9276$new_n2170;
    wire $abc$9276$new_n2171;
    wire $abc$9276$new_n2172;
    wire $abc$9276$new_n2173;
    wire $abc$9276$new_n2174;
    wire $abc$9276$new_n2175;
    wire $abc$9276$new_n2177;
    wire $abc$9276$new_n2178;
    wire $abc$9276$new_n2179;
    wire $abc$9276$new_n2180;
    wire $abc$9276$new_n2181;
    wire $abc$9276$new_n2182;
    wire $abc$9276$new_n2183;
    wire $abc$9276$new_n2184;
    wire $abc$9276$new_n2185;
    wire $abc$9276$new_n2186;
    wire $abc$9276$new_n2187;
    wire $abc$9276$new_n2188;
    wire $abc$9276$new_n2189;
    wire $abc$9276$new_n2190;
    wire $abc$9276$new_n2191;
    wire $abc$9276$new_n2192;
    wire $abc$9276$new_n2193;
    wire $abc$9276$new_n2194;
    wire $abc$9276$new_n2195;
    wire $abc$9276$new_n2196;
    wire $abc$9276$new_n2197;
    wire $abc$9276$new_n2198;
    wire $abc$9276$new_n2199;
    wire $abc$9276$new_n2200;
    wire $abc$9276$new_n2201;
    wire $abc$9276$new_n2202;
    wire $abc$9276$new_n2203;
    wire $abc$9276$new_n2204;
    wire $abc$9276$new_n2205;
    wire $abc$9276$new_n2206;
    wire $abc$9276$new_n2207;
    wire $abc$9276$new_n2208;
    wire $abc$9276$new_n2209;
    wire $abc$9276$new_n2210;
    wire $abc$9276$new_n2211;
    wire $abc$9276$new_n2212;
    wire $abc$9276$new_n2213;
    wire $abc$9276$new_n2214;
    wire $abc$9276$new_n2215;
    wire $abc$9276$new_n2216;
    wire $abc$9276$new_n2217;
    wire $abc$9276$new_n2218;
    wire $abc$9276$new_n2219;
    wire $abc$9276$new_n2220;
    wire $abc$9276$new_n2221;
    wire $abc$9276$new_n2222;
    wire $abc$9276$new_n2223;
    wire $abc$9276$new_n2224;
    wire $abc$9276$new_n2225;
    wire $abc$9276$new_n2226;
    wire $abc$9276$new_n2227;
    wire $abc$9276$new_n2228;
    wire $abc$9276$new_n2229;
    wire $abc$9276$new_n2230;
    wire $abc$9276$new_n2231;
    wire $abc$9276$new_n2232;
    wire $abc$9276$new_n2233;
    wire $abc$9276$new_n2234;
    wire $abc$9276$new_n2235;
    wire $abc$9276$new_n2236;
    wire $abc$9276$new_n2237;
    wire $abc$9276$new_n2238;
    wire $abc$9276$new_n2239;
    wire $abc$9276$new_n2240;
    wire $abc$9276$new_n2241;
    wire $abc$9276$new_n2242;
    wire $abc$9276$new_n2243;
    wire $abc$9276$new_n2244;
    wire $abc$9276$new_n2245;
    wire $abc$9276$new_n2246;
    wire $abc$9276$new_n2247;
    wire $abc$9276$new_n2248;
    wire $abc$9276$new_n2249;
    wire $abc$9276$new_n2250;
    wire $abc$9276$new_n2251;
    wire $abc$9276$new_n2252;
    wire $abc$9276$new_n2253;
    wire $abc$9276$new_n2254;
    wire $abc$9276$new_n2255;
    wire $abc$9276$new_n2256;
    wire $abc$9276$new_n2257;
    wire $abc$9276$new_n2258;
    wire $abc$9276$new_n2259;
    wire $abc$9276$new_n2260;
    wire $abc$9276$new_n2261;
    wire $abc$9276$new_n2262;
    wire $abc$9276$new_n2263;
    wire $abc$9276$new_n2264;
    wire $abc$9276$new_n2265;
    wire $abc$9276$new_n2266;
    wire $abc$9276$new_n2267;
    wire $abc$9276$new_n2268;
    wire $abc$9276$new_n2269;
    wire $abc$9276$new_n2270;
    wire $abc$9276$new_n2271;
    wire $abc$9276$new_n2272;
    wire $abc$9276$new_n2273;
    wire $abc$9276$new_n2274;
    wire $abc$9276$new_n2275;
    wire $abc$9276$new_n2276;
    wire $abc$9276$new_n2277;
    wire $abc$9276$new_n2278;
    wire $abc$9276$new_n2279;
    wire $abc$9276$new_n2280;
    wire $abc$9276$new_n2281;
    wire $abc$9276$new_n2282;
    wire $abc$9276$new_n2283;
    wire $abc$9276$new_n2284;
    wire $abc$9276$new_n2285;
    wire $abc$9276$new_n2286;
    wire $abc$9276$new_n2287;
    wire $abc$9276$new_n2288;
    wire $abc$9276$new_n2289;
    wire $abc$9276$new_n2290;
    wire $abc$9276$new_n2291;
    wire $abc$9276$new_n2292;
    wire $abc$9276$new_n2293;
    wire $abc$9276$new_n2294;
    wire $abc$9276$new_n2295;
    wire $abc$9276$new_n2296;
    wire $abc$9276$new_n2297;
    wire $abc$9276$new_n2298;
    wire $abc$9276$new_n2299;
    wire $abc$9276$new_n2300;
    wire $abc$9276$new_n2301;
    wire $abc$9276$new_n2302;
    wire $abc$9276$new_n2303;
    wire $abc$9276$new_n2304;
    wire $abc$9276$new_n2305;
    wire $abc$9276$new_n2307;
    wire $abc$9276$new_n2308;
    wire $abc$9276$new_n2309;
    wire $abc$9276$new_n2310;
    wire $abc$9276$new_n2311;
    wire $abc$9276$new_n2312;
    wire $abc$9276$new_n2313;
    wire $abc$9276$new_n2314;
    wire $abc$9276$new_n2315;
    wire $abc$9276$new_n2316;
    wire $abc$9276$new_n2317;
    wire $abc$9276$new_n2318;
    wire $abc$9276$new_n2319;
    wire $abc$9276$new_n2320;
    wire $abc$9276$new_n2321;
    wire $abc$9276$new_n2322;
    wire $abc$9276$new_n2323;
    wire $abc$9276$new_n2324;
    wire $abc$9276$new_n2325;
    wire $abc$9276$new_n2326;
    wire $abc$9276$new_n2327;
    wire $abc$9276$new_n2328;
    wire $abc$9276$new_n2329;
    wire $abc$9276$new_n2330;
    wire $abc$9276$new_n2331;
    wire $abc$9276$new_n2332;
    wire $abc$9276$new_n2333;
    wire $abc$9276$new_n2334;
    wire $abc$9276$new_n2335;
    wire $abc$9276$new_n2336;
    wire $abc$9276$new_n2337;
    wire $abc$9276$new_n2338;
    wire $abc$9276$new_n2339;
    wire $abc$9276$new_n2340;
    wire $abc$9276$new_n2341;
    wire $abc$9276$new_n2342;
    wire $abc$9276$new_n2343;
    wire $abc$9276$new_n2344;
    wire $abc$9276$new_n2345;
    wire $abc$9276$new_n2346;
    wire $abc$9276$new_n2347;
    wire $abc$9276$new_n2348;
    wire $abc$9276$new_n2349;
    wire $abc$9276$new_n2350;
    wire $abc$9276$new_n2351;
    wire $abc$9276$new_n2352;
    wire $abc$9276$new_n2353;
    wire $abc$9276$new_n2354;
    wire $abc$9276$new_n2355;
    wire $abc$9276$new_n2356;
    wire $abc$9276$new_n2357;
    wire $abc$9276$new_n2358;
    wire $abc$9276$new_n2359;
    wire $abc$9276$new_n2360;
    wire $abc$9276$new_n2361;
    wire $abc$9276$new_n2362;
    wire $abc$9276$new_n2363;
    wire $abc$9276$new_n2364;
    wire $abc$9276$new_n2365;
    wire $abc$9276$new_n2366;
    wire $abc$9276$new_n2367;
    wire $abc$9276$new_n2368;
    wire $abc$9276$new_n2369;
    wire $abc$9276$new_n2370;
    wire $abc$9276$new_n2371;
    wire $abc$9276$new_n2372;
    wire $abc$9276$new_n2373;
    wire $abc$9276$new_n2374;
    wire $abc$9276$new_n2375;
    wire $abc$9276$new_n2376;
    wire $abc$9276$new_n2377;
    wire $abc$9276$new_n2378;
    wire $abc$9276$new_n2379;
    wire $abc$9276$new_n2380;
    wire $abc$9276$new_n2381;
    wire $abc$9276$new_n2382;
    wire $abc$9276$new_n2383;
    wire $abc$9276$new_n2384;
    wire $abc$9276$new_n2385;
    wire $abc$9276$new_n2386;
    wire $abc$9276$new_n2387;
    wire $abc$9276$new_n2388;
    wire $abc$9276$new_n2389;
    wire $abc$9276$new_n2390;
    wire $abc$9276$new_n2391;
    wire $abc$9276$new_n2392;
    wire $abc$9276$new_n2393;
    wire $abc$9276$new_n2394;
    wire $abc$9276$new_n2395;
    wire $abc$9276$new_n2396;
    wire $abc$9276$new_n2397;
    wire $abc$9276$new_n2398;
    wire $abc$9276$new_n2399;
    wire $abc$9276$new_n2400;
    wire $abc$9276$new_n2401;
    wire $abc$9276$new_n2402;
    wire $abc$9276$new_n2403;
    wire $abc$9276$new_n2404;
    wire $abc$9276$new_n2405;
    wire $abc$9276$new_n2406;
    wire $abc$9276$new_n2407;
    wire $abc$9276$new_n2408;
    wire $abc$9276$new_n2409;
    wire $abc$9276$new_n2410;
    wire $abc$9276$new_n2411;
    wire $abc$9276$new_n2412;
    wire $abc$9276$new_n2413;
    wire $abc$9276$new_n2414;
    wire $abc$9276$new_n2415;
    wire $abc$9276$new_n2416;
    wire $abc$9276$new_n2417;
    wire $abc$9276$new_n2418;
    wire $abc$9276$new_n2419;
    wire $abc$9276$new_n2420;
    wire $abc$9276$new_n2421;
    wire $abc$9276$new_n2422;
    wire $abc$9276$new_n2423;
    wire $abc$9276$new_n2424;
    wire $abc$9276$new_n2425;
    wire $abc$9276$new_n2426;
    wire $abc$9276$new_n2427;
    wire $abc$9276$new_n2428;
    wire $abc$9276$new_n2429;
    wire $abc$9276$new_n2430;
    wire $abc$9276$new_n2431;
    wire $abc$9276$new_n2432;
    wire $abc$9276$new_n2433;
    wire $abc$9276$new_n2434;
    wire $abc$9276$new_n2435;
    wire $abc$9276$new_n2436;
    wire $abc$9276$new_n2437;
    wire $abc$9276$new_n2438;
    wire $abc$9276$new_n2439;
    wire $abc$9276$new_n2440;
    wire $abc$9276$new_n2441;
    wire $abc$9276$new_n2442;
    wire $abc$9276$new_n2443;
    wire $abc$9276$new_n2444;
    wire $abc$9276$new_n2445;
    wire $abc$9276$new_n2446;
    wire $abc$9276$new_n2447;
    wire $abc$9276$new_n2448;
    wire $abc$9276$new_n2449;
    wire $abc$9276$new_n2450;
    wire $abc$9276$new_n2451;
    wire $abc$9276$new_n2452;
    wire $abc$9276$new_n2453;
    wire $abc$9276$new_n2454;
    wire $abc$9276$new_n2455;
    wire $abc$9276$new_n2456;
    wire $abc$9276$new_n2457;
    wire $abc$9276$new_n2458;
    wire $abc$9276$new_n2459;
    wire $abc$9276$new_n2460;
    wire $abc$9276$new_n2461;
    wire $abc$9276$new_n2462;
    wire $abc$9276$new_n2463;
    wire $abc$9276$new_n2464;
    wire $abc$9276$new_n2465;
    wire $abc$9276$new_n2466;
    wire $abc$9276$new_n2467;
    wire $abc$9276$new_n2468;
    wire $abc$9276$new_n2469;
    wire $abc$9276$new_n2470;
    wire $abc$9276$new_n2471;
    wire $abc$9276$new_n2472;
    wire $abc$9276$new_n2473;
    wire $abc$9276$new_n2474;
    wire $abc$9276$new_n2475;
    wire $abc$9276$new_n2476;
    wire $abc$9276$new_n2477;
    wire $abc$9276$new_n2478;
    wire $abc$9276$new_n2479;
    wire $abc$9276$new_n2480;
    wire $abc$9276$new_n2481;
    wire $abc$9276$new_n2482;
    wire $abc$9276$new_n2483;
    wire $abc$9276$new_n2484;
    wire $abc$9276$new_n2485;
    wire $abc$9276$new_n2486;
    wire $abc$9276$new_n2487;
    wire $abc$9276$new_n2488;
    wire $abc$9276$new_n2489;
    wire $abc$9276$new_n2490;
    wire $abc$9276$new_n2491;
    wire $abc$9276$new_n2492;
    wire $abc$9276$new_n2493;
    wire $abc$9276$new_n2494;
    wire $abc$9276$new_n2495;
    wire $abc$9276$new_n2496;
    wire $abc$9276$new_n2497;
    wire $abc$9276$new_n2498;
    wire $abc$9276$new_n2499;
    wire $abc$9276$new_n2500;
    wire $abc$9276$new_n2501;
    wire $abc$9276$new_n2502;
    wire $abc$9276$new_n2503;
    wire $abc$9276$new_n2504;
    wire $abc$9276$new_n2505;
    wire $abc$9276$new_n2506;
    wire $abc$9276$new_n2507;
    wire $abc$9276$new_n2508;
    wire $abc$9276$new_n2509;
    wire $abc$9276$new_n2510;
    wire $abc$9276$new_n2511;
    wire $abc$9276$new_n2512;
    wire $abc$9276$new_n2513;
    wire $abc$9276$new_n2514;
    wire $abc$9276$new_n2515;
    wire $abc$9276$new_n2516;
    wire $abc$9276$new_n2517;
    wire $abc$9276$new_n2518;
    wire $abc$9276$new_n2519;
    wire $abc$9276$new_n2520;
    wire $abc$9276$new_n2521;
    wire $abc$9276$new_n2522;
    wire $abc$9276$new_n2523;
    wire $abc$9276$new_n2524;
    wire $abc$9276$new_n2525;
    wire $abc$9276$new_n2526;
    wire $abc$9276$new_n2527;
    wire $abc$9276$new_n2528;
    wire $abc$9276$new_n2529;
    wire $abc$9276$new_n2530;
    wire $abc$9276$new_n2531;
    wire $abc$9276$new_n2532;
    wire $abc$9276$new_n2533;
    wire $abc$9276$new_n2534;
    wire $abc$9276$new_n2535;
    wire $abc$9276$new_n2536;
    wire $abc$9276$new_n2537;
    wire $abc$9276$new_n2538;
    wire $abc$9276$new_n2539;
    wire $abc$9276$new_n2540;
    wire $abc$9276$new_n2541;
    wire $abc$9276$new_n2542;
    wire $abc$9276$new_n2543;
    wire $abc$9276$new_n2544;
    wire $abc$9276$new_n2545;
    wire $abc$9276$new_n2546;
    wire $abc$9276$new_n2547;
    wire $abc$9276$new_n2548;
    wire $abc$9276$new_n2549;
    wire $abc$9276$new_n2550;
    wire $abc$9276$new_n2551;
    wire $abc$9276$new_n2552;
    wire $abc$9276$new_n2553;
    wire $abc$9276$new_n2554;
    wire $abc$9276$new_n2555;
    wire $abc$9276$new_n2556;
    wire $abc$9276$new_n2557;
    wire $abc$9276$new_n2558;
    wire $abc$9276$new_n2559;
    wire $abc$9276$new_n2560;
    wire $abc$9276$new_n2561;
    wire $abc$9276$new_n2562;
    wire $abc$9276$new_n2563;
    wire $abc$9276$new_n2564;
    wire $abc$9276$new_n2565;
    wire $abc$9276$new_n2566;
    wire $abc$9276$new_n2567;
    wire $abc$9276$new_n2568;
    wire $abc$9276$new_n2569;
    wire $abc$9276$new_n2570;
    wire $abc$9276$new_n2571;
    wire $abc$9276$new_n2572;
    wire $abc$9276$new_n2573;
    wire $abc$9276$new_n2575;
    wire $abc$9276$new_n2576;
    wire $abc$9276$new_n2578;
    wire $abc$9276$new_n2579;
    wire $abc$9276$new_n2580;
    wire $abc$9276$new_n2581;
    wire $abc$9276$new_n2582;
    wire $abc$9276$new_n2584;
    wire $abc$9276$new_n2585;
    wire $abc$9276$new_n2586;
    wire $abc$9276$new_n2588;
    wire $abc$9276$new_n2589;
    wire $abc$9276$new_n2590;
    wire $abc$9276$new_n2592;
    wire $abc$9276$new_n2593;
    wire $abc$9276$new_n2594;
    wire $abc$9276$new_n2596;
    wire $abc$9276$new_n2597;
    wire $abc$9276$new_n2598;
    wire $abc$9276$new_n2599;
    wire $abc$9276$new_n2600;
    wire $abc$9276$new_n2602;
    wire $abc$9276$new_n2603;
    wire $abc$9276$new_n2604;
    wire $abc$9276$new_n2605;
    wire $abc$9276$new_n2606;
    wire $abc$9276$new_n2608;
    wire $abc$9276$new_n2609;
    wire $abc$9276$new_n2610;
    wire $abc$9276$new_n2611;
    wire $abc$9276$new_n2612;
    wire $abc$9276$new_n2614;
    wire $abc$9276$new_n2615;
    wire $abc$9276$new_n2617;
    wire $abc$9276$new_n2618;
    wire $abc$9276$new_n2619;
    wire $abc$9276$new_n2620;
    wire $abc$9276$new_n2621;
    wire $abc$9276$new_n2622;
    wire $abc$9276$new_n2623;
    wire $abc$9276$new_n2624;
    wire $abc$9276$new_n2625;
    wire $abc$9276$new_n2626;
    wire $abc$9276$new_n2627;
    wire $abc$9276$new_n2628;
    wire $abc$9276$new_n2629;
    wire $abc$9276$new_n2630;
    wire $abc$9276$new_n2631;
    wire $abc$9276$new_n2633;
    wire $abc$9276$new_n2634;
    wire $abc$9276$new_n2635;
    wire $abc$9276$new_n2636;
    wire $abc$9276$new_n2637;
    wire $abc$9276$new_n2638;
    wire $abc$9276$new_n2640;
    wire $abc$9276$new_n2641;
    wire $abc$9276$new_n2642;
    wire $abc$9276$new_n2643;
    wire $abc$9276$new_n2645;
    wire $abc$9276$new_n2646;
    wire $abc$9276$new_n2647;
    wire $abc$9276$new_n2648;
    wire $abc$9276$new_n2649;
    wire $abc$9276$new_n2650;
    wire $abc$9276$new_n2651;
    wire $abc$9276$new_n2652;
    wire $abc$9276$new_n2654;
    wire $abc$9276$new_n2655;
    wire $abc$9276$new_n2656;
    wire $abc$9276$new_n2657;
    wire $abc$9276$new_n2658;
    wire $abc$9276$new_n2659;
    wire $abc$9276$new_n2660;
    wire $abc$9276$new_n2661;
    wire $abc$9276$new_n2662;
    wire $abc$9276$new_n2663;
    wire $abc$9276$new_n2664;
    wire $abc$9276$new_n2665;
    wire $abc$9276$new_n2666;
    wire $abc$9276$new_n2667;
    wire $abc$9276$new_n2668;
    wire $abc$9276$new_n2669;
    wire $abc$9276$new_n2671;
    wire $abc$9276$new_n2672;
    wire $abc$9276$new_n2673;
    wire $abc$9276$new_n2674;
    wire $abc$9276$new_n2675;
    wire $abc$9276$new_n2676;
    wire $abc$9276$new_n2678;
    wire $abc$9276$new_n2679;
    wire $abc$9276$new_n2680;
    wire $abc$9276$new_n2681;
    wire $abc$9276$new_n2682;
    wire $abc$9276$new_n2683;
    wire $abc$9276$new_n2684;
    wire $abc$9276$new_n2685;
    wire $abc$9276$new_n2686;
    wire $abc$9276$new_n2687;
    wire $abc$9276$new_n2688;
    wire $abc$9276$new_n2689;
    wire $abc$9276$new_n2690;
    wire $abc$9276$new_n2691;
    wire $abc$9276$new_n2693;
    wire $abc$9276$new_n2694;
    wire $abc$9276$new_n2695;
    wire $abc$9276$new_n2696;
    wire $abc$9276$new_n2697;
    wire $abc$9276$new_n2698;
    wire $abc$9276$new_n2699;
    wire $abc$9276$new_n2700;
    wire $abc$9276$new_n2701;
    wire $abc$9276$new_n2702;
    wire $abc$9276$new_n2703;
    wire $abc$9276$new_n2705;
    wire $abc$9276$new_n2706;
    wire $abc$9276$new_n2707;
    wire $abc$9276$new_n2708;
    wire $abc$9276$new_n2709;
    wire $abc$9276$new_n2710;
    wire $abc$9276$new_n2711;
    wire $abc$9276$new_n2712;
    wire $abc$9276$new_n2713;
    wire $abc$9276$new_n2714;
    wire $abc$9276$new_n2715;
    wire $abc$9276$new_n2717;
    wire $abc$9276$new_n2718;
    wire $abc$9276$new_n2719;
    wire $abc$9276$new_n2720;
    wire $abc$9276$new_n2721;
    wire $abc$9276$new_n2722;
    wire $abc$9276$new_n2723;
    wire $abc$9276$new_n2724;
    wire $abc$9276$new_n2725;
    wire $abc$9276$new_n2727;
    wire $abc$9276$new_n2728;
    wire $abc$9276$new_n2729;
    wire $abc$9276$new_n2730;
    wire $abc$9276$new_n2731;
    wire $abc$9276$new_n2732;
    wire $abc$9276$new_n2733;
    wire $abc$9276$new_n2734;
    wire $abc$9276$new_n2735;
    wire $abc$9276$new_n2736;
    wire $abc$9276$new_n2737;
    wire $abc$9276$new_n2738;
    wire $abc$9276$new_n2740;
    wire $abc$9276$new_n2741;
    wire $abc$9276$new_n2742;
    wire $abc$9276$new_n2743;
    wire $abc$9276$new_n2744;
    wire $abc$9276$new_n2745;
    wire $abc$9276$new_n2746;
    wire $abc$9276$new_n2747;
    wire $abc$9276$new_n2748;
    wire $abc$9276$new_n2749;
    wire $abc$9276$new_n2751;
    wire $abc$9276$new_n2752;
    wire $abc$9276$new_n2753;
    wire $abc$9276$new_n2754;
    wire $abc$9276$new_n2755;
    wire $abc$9276$new_n2756;
    wire $abc$9276$new_n2757;
    wire $abc$9276$new_n2758;
    wire $abc$9276$new_n2759;
    wire $abc$9276$new_n2760;
    wire $abc$9276$new_n2761;
    wire $abc$9276$new_n2763;
    wire $abc$9276$new_n2764;
    wire $abc$9276$new_n2765;
    wire $abc$9276$new_n2766;
    wire $abc$9276$new_n2767;
    wire $abc$9276$new_n2768;
    wire $abc$9276$new_n2769;
    wire $abc$9276$new_n2770;
    wire $abc$9276$new_n2771;
    wire $abc$9276$new_n2772;
    wire $abc$9276$new_n2773;
    wire $abc$9276$new_n2775;
    wire $abc$9276$new_n346;
    wire $abc$9276$new_n347;
    wire $abc$9276$new_n348;
    wire $abc$9276$new_n349;
    wire $abc$9276$new_n350;
    wire $abc$9276$new_n351;
    wire $abc$9276$new_n352;
    wire $abc$9276$new_n353;
    wire $abc$9276$new_n354;
    wire $abc$9276$new_n355;
    wire $abc$9276$new_n356;
    wire $abc$9276$new_n357;
    wire $abc$9276$new_n358;
    wire $abc$9276$new_n359;
    wire $abc$9276$new_n360;
    wire $abc$9276$new_n361;
    wire $abc$9276$new_n362;
    wire $abc$9276$new_n363;
    wire $abc$9276$new_n364;
    wire $abc$9276$new_n365;
    wire $abc$9276$new_n366;
    wire $abc$9276$new_n367;
    wire $abc$9276$new_n368;
    wire $abc$9276$new_n369;
    wire $abc$9276$new_n370;
    wire $abc$9276$new_n371;
    wire $abc$9276$new_n372;
    wire $abc$9276$new_n373;
    wire $abc$9276$new_n374;
    wire $abc$9276$new_n375;
    wire $abc$9276$new_n376;
    wire $abc$9276$new_n377;
    wire $abc$9276$new_n378;
    wire $abc$9276$new_n379;
    wire $abc$9276$new_n380;
    wire $abc$9276$new_n381;
    wire $abc$9276$new_n382;
    wire $abc$9276$new_n383;
    wire $abc$9276$new_n384;
    wire $abc$9276$new_n385;
    wire $abc$9276$new_n386;
    wire $abc$9276$new_n387;
    wire $abc$9276$new_n388;
    wire $abc$9276$new_n389;
    wire $abc$9276$new_n390;
    wire $abc$9276$new_n391;
    wire $abc$9276$new_n392;
    wire $abc$9276$new_n393;
    wire $abc$9276$new_n394;
    wire $abc$9276$new_n395;
    wire $abc$9276$new_n396;
    wire $abc$9276$new_n397;
    wire $abc$9276$new_n398;
    wire $abc$9276$new_n399;
    wire $abc$9276$new_n400;
    wire $abc$9276$new_n401;
    wire $abc$9276$new_n402;
    wire $abc$9276$new_n403;
    wire $abc$9276$new_n404;
    wire $abc$9276$new_n405;
    wire $abc$9276$new_n406;
    wire $abc$9276$new_n407;
    wire $abc$9276$new_n408;
    wire $abc$9276$new_n409;
    wire $abc$9276$new_n410;
    wire $abc$9276$new_n411;
    wire $abc$9276$new_n412;
    wire $abc$9276$new_n413;
    wire $abc$9276$new_n414;
    wire $abc$9276$new_n415;
    wire $abc$9276$new_n416;
    wire $abc$9276$new_n417;
    wire $abc$9276$new_n418;
    wire $abc$9276$new_n419;
    wire $abc$9276$new_n420;
    wire $abc$9276$new_n421;
    wire $abc$9276$new_n422;
    wire $abc$9276$new_n423;
    wire $abc$9276$new_n424;
    wire $abc$9276$new_n425;
    wire $abc$9276$new_n426;
    wire $abc$9276$new_n427;
    wire $abc$9276$new_n428;
    wire $abc$9276$new_n429;
    wire $abc$9276$new_n430;
    wire $abc$9276$new_n431;
    wire $abc$9276$new_n432;
    wire $abc$9276$new_n433;
    wire $abc$9276$new_n434;
    wire $abc$9276$new_n435;
    wire $abc$9276$new_n436;
    wire $abc$9276$new_n437;
    wire $abc$9276$new_n438;
    wire $abc$9276$new_n439;
    wire $abc$9276$new_n440;
    wire $abc$9276$new_n441;
    wire $abc$9276$new_n442;
    wire $abc$9276$new_n443;
    wire $abc$9276$new_n444;
    wire $abc$9276$new_n445;
    wire $abc$9276$new_n446;
    wire $abc$9276$new_n447;
    wire $abc$9276$new_n448;
    wire $abc$9276$new_n449;
    wire $abc$9276$new_n450;
    wire $abc$9276$new_n451;
    wire $abc$9276$new_n452;
    wire $abc$9276$new_n453;
    wire $abc$9276$new_n454;
    wire $abc$9276$new_n455;
    wire $abc$9276$new_n456;
    wire $abc$9276$new_n457;
    wire $abc$9276$new_n458;
    wire $abc$9276$new_n459;
    wire $abc$9276$new_n460;
    wire $abc$9276$new_n461;
    wire $abc$9276$new_n462;
    wire $abc$9276$new_n463;
    wire $abc$9276$new_n464;
    wire $abc$9276$new_n465;
    wire $abc$9276$new_n466;
    wire $abc$9276$new_n467;
    wire $abc$9276$new_n468;
    wire $abc$9276$new_n469;
    wire $abc$9276$new_n470;
    wire $abc$9276$new_n471;
    wire $abc$9276$new_n472;
    wire $abc$9276$new_n473;
    wire $abc$9276$new_n474;
    wire $abc$9276$new_n475;
    wire $abc$9276$new_n476;
    wire $abc$9276$new_n477;
    wire $abc$9276$new_n478;
    wire $abc$9276$new_n479;
    wire $abc$9276$new_n480;
    wire $abc$9276$new_n481;
    wire $abc$9276$new_n482;
    wire $abc$9276$new_n483;
    wire $abc$9276$new_n484;
    wire $abc$9276$new_n485;
    wire $abc$9276$new_n486;
    wire $abc$9276$new_n487;
    wire $abc$9276$new_n489;
    wire $abc$9276$new_n490;
    wire $abc$9276$new_n491;
    wire $abc$9276$new_n492;
    wire $abc$9276$new_n493;
    wire $abc$9276$new_n494;
    wire $abc$9276$new_n496;
    wire $abc$9276$new_n497;
    wire $abc$9276$new_n498;
    wire $abc$9276$new_n499;
    wire $abc$9276$new_n500;
    wire $abc$9276$new_n501;
    wire $abc$9276$new_n502;
    wire $abc$9276$new_n503;
    wire $abc$9276$new_n504;
    wire $abc$9276$new_n505;
    wire $abc$9276$new_n507;
    wire $abc$9276$new_n508;
    wire $abc$9276$new_n509;
    wire $abc$9276$new_n510;
    wire $abc$9276$new_n511;
    wire $abc$9276$new_n512;
    wire $abc$9276$new_n514;
    wire $abc$9276$new_n515;
    wire $abc$9276$new_n516;
    wire $abc$9276$new_n517;
    wire $abc$9276$new_n518;
    wire $abc$9276$new_n519;
    wire $abc$9276$new_n520;
    wire $abc$9276$new_n521;
    wire $abc$9276$new_n522;
    wire $abc$9276$new_n523;
    wire $abc$9276$new_n524;
    wire $abc$9276$new_n525;
    wire $abc$9276$new_n527;
    wire $abc$9276$new_n528;
    wire $abc$9276$new_n529;
    wire $abc$9276$new_n530;
    wire $abc$9276$new_n531;
    wire $abc$9276$new_n532;
    wire $abc$9276$new_n534;
    wire $abc$9276$new_n535;
    wire $abc$9276$new_n536;
    wire $abc$9276$new_n537;
    wire $abc$9276$new_n538;
    wire $abc$9276$new_n539;
    wire $abc$9276$new_n540;
    wire $abc$9276$new_n541;
    wire $abc$9276$new_n542;
    wire $abc$9276$new_n543;
    wire $abc$9276$new_n544;
    wire $abc$9276$new_n545;
    wire $abc$9276$new_n547;
    wire $abc$9276$new_n548;
    wire $abc$9276$new_n549;
    wire $abc$9276$new_n550;
    wire $abc$9276$new_n551;
    wire $abc$9276$new_n552;
    wire $abc$9276$new_n554;
    wire $abc$9276$new_n555;
    wire $abc$9276$new_n556;
    wire $abc$9276$new_n557;
    wire $abc$9276$new_n558;
    wire $abc$9276$new_n559;
    wire $abc$9276$new_n560;
    wire $abc$9276$new_n561;
    wire $abc$9276$new_n562;
    wire $abc$9276$new_n563;
    wire $abc$9276$new_n564;
    wire $abc$9276$new_n565;
    wire $abc$9276$new_n566;
    wire $abc$9276$new_n567;
    wire $abc$9276$new_n568;
    wire $abc$9276$new_n570;
    wire $abc$9276$new_n571;
    wire $abc$9276$new_n572;
    wire $abc$9276$new_n573;
    wire $abc$9276$new_n574;
    wire $abc$9276$new_n575;
    wire $abc$9276$new_n577;
    wire $abc$9276$new_n578;
    wire $abc$9276$new_n579;
    wire $abc$9276$new_n580;
    wire $abc$9276$new_n581;
    wire $abc$9276$new_n582;
    wire $abc$9276$new_n583;
    wire $abc$9276$new_n584;
    wire $abc$9276$new_n585;
    wire $abc$9276$new_n586;
    wire $abc$9276$new_n588;
    wire $abc$9276$new_n589;
    wire $abc$9276$new_n590;
    wire $abc$9276$new_n591;
    wire $abc$9276$new_n592;
    wire $abc$9276$new_n593;
    wire $abc$9276$new_n595;
    wire $abc$9276$new_n596;
    wire $abc$9276$new_n597;
    wire $abc$9276$new_n598;
    wire $abc$9276$new_n599;
    wire $abc$9276$new_n600;
    wire $abc$9276$new_n601;
    wire $abc$9276$new_n602;
    wire $abc$9276$new_n603;
    wire $abc$9276$new_n604;
    wire $abc$9276$new_n605;
    wire $abc$9276$new_n606;
    wire $abc$9276$new_n608;
    wire $abc$9276$new_n609;
    wire $abc$9276$new_n610;
    wire $abc$9276$new_n611;
    wire $abc$9276$new_n612;
    wire $abc$9276$new_n613;
    wire $abc$9276$new_n615;
    wire $abc$9276$new_n616;
    wire $abc$9276$new_n617;
    wire $abc$9276$new_n618;
    wire $abc$9276$new_n619;
    wire $abc$9276$new_n620;
    wire $abc$9276$new_n621;
    wire $abc$9276$new_n622;
    wire $abc$9276$new_n623;
    wire $abc$9276$new_n624;
    wire $abc$9276$new_n626;
    wire $abc$9276$new_n627;
    wire $abc$9276$new_n628;
    wire $abc$9276$new_n629;
    wire $abc$9276$new_n630;
    wire $abc$9276$new_n631;
    wire $abc$9276$new_n633;
    wire $abc$9276$new_n634;
    wire $abc$9276$new_n635;
    wire $abc$9276$new_n637;
    wire $abc$9276$new_n638;
    wire $abc$9276$new_n640;
    wire $abc$9276$new_n641;
    wire $abc$9276$new_n643;
    wire $abc$9276$new_n644;
    wire $abc$9276$new_n646;
    wire $abc$9276$new_n647;
    wire $abc$9276$new_n649;
    wire $abc$9276$new_n650;
    wire $abc$9276$new_n652;
    wire $abc$9276$new_n653;
    wire $abc$9276$new_n655;
    wire $abc$9276$new_n656;
    wire $abc$9276$new_n658;
    wire $abc$9276$new_n659;
    wire $abc$9276$new_n660;
    wire $abc$9276$new_n661;
    wire $abc$9276$new_n663;
    wire $abc$9276$new_n664;
    wire $abc$9276$new_n666;
    wire $abc$9276$new_n667;
    wire $abc$9276$new_n669;
    wire $abc$9276$new_n670;
    wire $abc$9276$new_n672;
    wire $abc$9276$new_n673;
    wire $abc$9276$new_n675;
    wire $abc$9276$new_n676;
    wire $abc$9276$new_n678;
    wire $abc$9276$new_n679;
    wire $abc$9276$new_n681;
    wire $abc$9276$new_n682;
    wire $abc$9276$new_n684;
    wire $abc$9276$new_n685;
    wire $abc$9276$new_n686;
    wire $abc$9276$new_n687;
    wire $abc$9276$new_n689;
    wire $abc$9276$new_n690;
    wire $abc$9276$new_n692;
    wire $abc$9276$new_n693;
    wire $abc$9276$new_n695;
    wire $abc$9276$new_n696;
    wire $abc$9276$new_n698;
    wire $abc$9276$new_n699;
    wire $abc$9276$new_n701;
    wire $abc$9276$new_n702;
    wire $abc$9276$new_n704;
    wire $abc$9276$new_n705;
    wire $abc$9276$new_n707;
    wire $abc$9276$new_n708;
    wire $abc$9276$new_n710;
    wire $abc$9276$new_n711;
    wire $abc$9276$new_n712;
    wire $abc$9276$new_n713;
    wire $abc$9276$new_n714;
    wire $abc$9276$new_n715;
    wire $abc$9276$new_n716;
    wire $abc$9276$new_n717;
    wire $abc$9276$new_n718;
    wire $abc$9276$new_n719;
    wire $abc$9276$new_n720;
    wire $abc$9276$new_n721;
    wire $abc$9276$new_n722;
    wire $abc$9276$new_n723;
    wire $abc$9276$new_n724;
    wire $abc$9276$new_n725;
    wire $abc$9276$new_n726;
    wire $abc$9276$new_n727;
    wire $abc$9276$new_n728;
    wire $abc$9276$new_n729;
    wire $abc$9276$new_n730;
    wire $abc$9276$new_n731;
    wire $abc$9276$new_n732;
    wire $abc$9276$new_n733;
    wire $abc$9276$new_n734;
    wire $abc$9276$new_n735;
    wire $abc$9276$new_n736;
    wire $abc$9276$new_n737;
    wire $abc$9276$new_n738;
    wire $abc$9276$new_n739;
    wire $abc$9276$new_n740;
    wire $abc$9276$new_n741;
    wire $abc$9276$new_n742;
    wire $abc$9276$new_n743;
    wire $abc$9276$new_n744;
    wire $abc$9276$new_n745;
    wire $abc$9276$new_n746;
    wire $abc$9276$new_n747;
    wire $abc$9276$new_n748;
    wire $abc$9276$new_n749;
    wire $abc$9276$new_n750;
    wire $abc$9276$new_n752;
    wire $abc$9276$new_n753;
    wire $abc$9276$new_n754;
    wire $abc$9276$new_n755;
    wire $abc$9276$new_n756;
    wire $abc$9276$new_n757;
    wire $abc$9276$new_n758;
    wire $abc$9276$new_n759;
    wire $abc$9276$new_n760;
    wire $abc$9276$new_n761;
    wire $abc$9276$new_n762;
    wire $abc$9276$new_n763;
    wire $abc$9276$new_n764;
    wire $abc$9276$new_n765;
    wire $abc$9276$new_n766;
    wire $abc$9276$new_n767;
    wire $abc$9276$new_n768;
    wire $abc$9276$new_n769;
    wire $abc$9276$new_n770;
    wire $abc$9276$new_n771;
    wire $abc$9276$new_n772;
    wire $abc$9276$new_n773;
    wire $abc$9276$new_n774;
    wire $abc$9276$new_n775;
    wire $abc$9276$new_n776;
    wire $abc$9276$new_n777;
    wire $abc$9276$new_n778;
    wire $abc$9276$new_n779;
    wire $abc$9276$new_n780;
    wire $abc$9276$new_n781;
    wire $abc$9276$new_n782;
    wire $abc$9276$new_n783;
    wire $abc$9276$new_n784;
    wire $abc$9276$new_n785;
    wire $abc$9276$new_n786;
    wire $abc$9276$new_n787;
    wire $abc$9276$new_n788;
    wire $abc$9276$new_n789;
    wire $abc$9276$new_n790;
    wire $abc$9276$new_n791;
    wire $abc$9276$new_n792;
    wire $abc$9276$new_n793;
    wire $abc$9276$new_n794;
    wire $abc$9276$new_n795;
    wire $abc$9276$new_n796;
    wire $abc$9276$new_n797;
    wire $abc$9276$new_n798;
    wire $abc$9276$new_n799;
    wire $abc$9276$new_n800;
    wire $abc$9276$new_n801;
    wire $abc$9276$new_n802;
    wire $abc$9276$new_n803;
    wire $abc$9276$new_n804;
    wire $abc$9276$new_n805;
    wire $abc$9276$new_n806;
    wire $abc$9276$new_n807;
    wire $abc$9276$new_n808;
    wire $abc$9276$new_n809;
    wire $abc$9276$new_n810;
    wire $abc$9276$new_n811;
    wire $abc$9276$new_n812;
    wire $abc$9276$new_n813;
    wire $abc$9276$new_n814;
    wire $abc$9276$new_n815;
    wire $abc$9276$new_n816;
    wire $abc$9276$new_n817;
    wire $abc$9276$new_n818;
    wire $abc$9276$new_n820;
    wire $abc$9276$new_n821;
    wire $abc$9276$new_n822;
    wire $abc$9276$new_n823;
    wire $abc$9276$new_n825;
    wire $abc$9276$new_n826;
    wire $abc$9276$new_n827;
    wire $abc$9276$new_n828;
    wire $abc$9276$new_n829;
    wire $abc$9276$new_n830;
    wire $abc$9276$new_n831;
    wire $abc$9276$new_n833;
    wire $abc$9276$new_n834;
    wire $abc$9276$new_n835;
    wire $abc$9276$new_n836;
    wire $abc$9276$new_n838;
    wire $abc$9276$new_n839;
    wire $abc$9276$new_n840;
    wire $abc$9276$new_n842;
    wire $abc$9276$new_n843;
    wire $abc$9276$new_n845;
    wire $abc$9276$new_n846;
    wire $abc$9276$new_n847;
    wire $abc$9276$new_n849;
    wire $abc$9276$new_n850;
    wire $abc$9276$new_n852;
    wire $abc$9276$new_n853;
    wire $abc$9276$new_n854;
    wire $abc$9276$new_n855;
    wire $abc$9276$new_n857;
    wire $abc$9276$new_n858;
    wire $abc$9276$new_n859;
    wire $abc$9276$new_n860;
    wire $abc$9276$new_n861;
    wire $abc$9276$new_n863;
    wire $abc$9276$new_n864;
    wire $abc$9276$new_n865;
    wire $abc$9276$new_n866;
    wire $abc$9276$new_n867;
    wire $abc$9276$new_n868;
    wire $abc$9276$new_n869;
    wire $abc$9276$new_n870;
    wire $abc$9276$new_n871;
    wire $abc$9276$new_n872;
    wire $abc$9276$new_n874;
    wire $abc$9276$new_n875;
    wire $abc$9276$new_n876;
    wire $abc$9276$new_n878;
    wire $abc$9276$new_n879;
    wire $abc$9276$new_n880;
    wire $abc$9276$new_n881;
    wire $abc$9276$new_n882;
    wire $abc$9276$new_n883;
    wire $abc$9276$new_n884;
    wire $abc$9276$new_n885;
    wire $abc$9276$new_n886;
    wire $abc$9276$new_n887;
    wire $abc$9276$new_n888;
    wire $abc$9276$new_n889;
    wire $abc$9276$new_n890;
    wire $abc$9276$new_n891;
    wire $abc$9276$new_n892;
    wire $abc$9276$new_n893;
    wire $abc$9276$new_n894;
    wire $abc$9276$new_n895;
    wire $abc$9276$new_n896;
    wire $abc$9276$new_n898;
    wire $abc$9276$new_n900;
    wire $abc$9276$new_n901;
    wire $abc$9276$new_n902;
    wire $abc$9276$new_n903;
    wire $abc$9276$new_n904;
    wire $abc$9276$new_n905;
    wire $abc$9276$new_n907;
    wire $abc$9276$new_n908;
    wire $abc$9276$new_n909;
    wire $abc$9276$new_n911;
    wire $abc$9276$new_n912;
    wire $abc$9276$new_n913;
    wire $abc$9276$new_n914;
    wire $abc$9276$new_n915;
    wire $abc$9276$new_n916;
    wire $abc$9276$new_n918;
    wire $abc$9276$new_n919;
    wire $abc$9276$new_n920;
    wire $abc$9276$new_n922;
    wire $abc$9276$new_n923;
    wire $abc$9276$new_n924;
    wire $abc$9276$new_n926;
    wire $abc$9276$new_n927;
    wire $abc$9276$new_n928;
    wire $abc$9276$new_n929;
    wire $abc$9276$new_n930;
    wire $abc$9276$new_n932;
    wire $abc$9276$new_n933;
    wire $abc$9276$new_n934;
    wire $abc$9276$new_n935;
    wire $abc$9276$new_n936;
    wire $abc$9276$new_n937;
    wire $abc$9276$new_n938;
    wire $abc$9276$new_n939;
    wire $abc$9276$new_n940;
    wire $abc$9276$new_n941;
    wire $abc$9276$new_n942;
    wire $abc$9276$new_n943;
    wire $abc$9276$new_n944;
    wire $abc$9276$new_n946;
    wire $abc$9276$new_n947;
    wire $abc$9276$new_n948;
    wire $abc$9276$new_n949;
    wire $abc$9276$new_n950;
    wire $abc$9276$new_n951;
    wire $abc$9276$new_n952;
    wire $abc$9276$new_n953;
    wire $abc$9276$new_n954;
    wire $abc$9276$new_n955;
    wire $abc$9276$new_n956;
    wire $abc$9276$new_n957;
    wire $abc$9276$new_n958;
    wire $abc$9276$new_n959;
    wire $abc$9276$new_n960;
    wire $abc$9276$new_n961;
    wire $abc$9276$new_n962;
    wire $abc$9276$new_n963;
    wire $abc$9276$new_n964;
    wire $abc$9276$new_n965;
    wire $abc$9276$new_n966;
    wire $abc$9276$new_n967;
    wire $abc$9276$new_n968;
    wire $abc$9276$new_n969;
    wire $abc$9276$new_n970;
    wire $abc$9276$new_n971;
    wire $abc$9276$new_n972;
    wire $abc$9276$new_n973;
    wire $abc$9276$new_n975;
    wire $abc$9276$new_n976;
    wire $abc$9276$new_n977;
    wire $abc$9276$new_n978;
    wire $abc$9276$new_n979;
    wire $abc$9276$new_n980;
    wire $abc$9276$new_n981;
    wire $abc$9276$new_n982;
    wire $abc$9276$new_n983;
    wire $abc$9276$new_n984;
    wire $abc$9276$new_n985;
    wire $abc$9276$new_n986;
    wire $abc$9276$new_n987;
    wire $abc$9276$new_n988;
    wire $abc$9276$new_n989;
    wire $abc$9276$new_n990;
    wire $abc$9276$new_n991;
    wire $abc$9276$new_n992;
    wire $abc$9276$new_n993;
    wire $abc$9276$new_n994;
    wire $abc$9276$new_n995;
    wire $abc$9276$new_n996;
    wire $abc$9276$new_n997;
    wire $abc$9276$new_n998;
    wire $abc$9276$new_n999;
    wire $auto$dfflibmap.cc:532:dfflibmap$9112;
    wire $auto$dfflibmap.cc:532:dfflibmap$9113;
    wire $auto$dfflibmap.cc:532:dfflibmap$9114;
    wire $auto$dfflibmap.cc:532:dfflibmap$9115;
    wire $auto$dfflibmap.cc:532:dfflibmap$9116;
    wire $auto$dfflibmap.cc:532:dfflibmap$9117;
    wire $auto$dfflibmap.cc:532:dfflibmap$9118;
    wire $auto$dfflibmap.cc:532:dfflibmap$9119;
    wire $auto$dfflibmap.cc:532:dfflibmap$9122;
    wire $auto$dfflibmap.cc:532:dfflibmap$9123;
    wire $auto$dfflibmap.cc:532:dfflibmap$9124;
    wire $auto$dfflibmap.cc:532:dfflibmap$9125;
    wire $auto$dfflibmap.cc:532:dfflibmap$9126;
    wire $auto$dfflibmap.cc:532:dfflibmap$9127;
    wire $auto$dfflibmap.cc:532:dfflibmap$9128;
    wire $auto$dfflibmap.cc:532:dfflibmap$9129;
    wire $auto$dfflibmap.cc:532:dfflibmap$9130;
    wire $auto$dfflibmap.cc:532:dfflibmap$9131;
    wire $auto$dfflibmap.cc:532:dfflibmap$9144;
    wire $auto$dfflibmap.cc:532:dfflibmap$9145;
    wire $auto$dfflibmap.cc:532:dfflibmap$9146;
    wire $auto$dfflibmap.cc:532:dfflibmap$9147;
    wire $auto$dfflibmap.cc:532:dfflibmap$9148;
    wire $auto$dfflibmap.cc:532:dfflibmap$9149;
    wire $auto$dfflibmap.cc:532:dfflibmap$9150;
    wire $auto$dfflibmap.cc:532:dfflibmap$9151;
    wire $auto$dfflibmap.cc:532:dfflibmap$9152;
    wire $auto$dfflibmap.cc:532:dfflibmap$9153;
    wire $auto$dfflibmap.cc:532:dfflibmap$9154;
    wire $auto$dfflibmap.cc:532:dfflibmap$9155;
    wire $auto$dfflibmap.cc:532:dfflibmap$9156;
    wire $auto$dfflibmap.cc:532:dfflibmap$9157;
    wire $auto$dfflibmap.cc:532:dfflibmap$9158;
    wire $auto$dfflibmap.cc:532:dfflibmap$9159;
    wire $auto$dfflibmap.cc:532:dfflibmap$9162;
    wire $auto$dfflibmap.cc:532:dfflibmap$9163;
    wire $auto$dfflibmap.cc:532:dfflibmap$9164;
    wire $auto$dfflibmap.cc:532:dfflibmap$9165;
    wire $auto$dfflibmap.cc:532:dfflibmap$9166;
    wire $auto$dfflibmap.cc:532:dfflibmap$9167;
    wire $auto$dfflibmap.cc:532:dfflibmap$9168;
    wire $auto$dfflibmap.cc:532:dfflibmap$9169;
    wire $auto$dfflibmap.cc:532:dfflibmap$9178;
    wire $auto$dfflibmap.cc:532:dfflibmap$9179;
    wire $auto$dfflibmap.cc:532:dfflibmap$9186;
    wire $auto$dfflibmap.cc:532:dfflibmap$9187;
    wire $auto$dfflibmap.cc:532:dfflibmap$9188;
    wire $auto$dfflibmap.cc:532:dfflibmap$9189;
    wire $auto$dfflibmap.cc:532:dfflibmap$9190;
    wire $auto$dfflibmap.cc:532:dfflibmap$9191;
    wire $auto$dfflibmap.cc:532:dfflibmap$9192;
    wire $auto$dfflibmap.cc:532:dfflibmap$9193;
    wire $auto$dfflibmap.cc:532:dfflibmap$9194;
    wire $auto$dfflibmap.cc:532:dfflibmap$9195;
    wire $auto$dfflibmap.cc:532:dfflibmap$9196;
    wire $auto$dfflibmap.cc:532:dfflibmap$9197;
    wire $auto$dfflibmap.cc:532:dfflibmap$9198;
    wire $auto$dfflibmap.cc:532:dfflibmap$9199;
    wire $auto$dfflibmap.cc:532:dfflibmap$9200;
    wire $auto$dfflibmap.cc:532:dfflibmap$9201;
    wire $auto$dfflibmap.cc:532:dfflibmap$9202;
    wire $auto$dfflibmap.cc:532:dfflibmap$9203;
    wire $auto$dfflibmap.cc:532:dfflibmap$9204;
    wire $auto$dfflibmap.cc:532:dfflibmap$9205;
    wire $auto$dfflibmap.cc:532:dfflibmap$9208;
    wire $auto$dfflibmap.cc:532:dfflibmap$9209;
    wire $auto$dfflibmap.cc:532:dfflibmap$9212;
    wire $auto$dfflibmap.cc:532:dfflibmap$9213;
    wire $auto$dfflibmap.cc:532:dfflibmap$9214;
    wire $auto$dfflibmap.cc:532:dfflibmap$9215;
    wire $auto$dfflibmap.cc:532:dfflibmap$9216;
    wire $auto$dfflibmap.cc:532:dfflibmap$9217;
    wire $auto$dfflibmap.cc:532:dfflibmap$9218;
    wire $auto$dfflibmap.cc:532:dfflibmap$9219;
    wire $auto$dfflibmap.cc:532:dfflibmap$9220;
    wire $auto$dfflibmap.cc:532:dfflibmap$9221;
    wire $auto$dfflibmap.cc:532:dfflibmap$9222;
    wire $auto$dfflibmap.cc:532:dfflibmap$9223;
    wire $auto$dfflibmap.cc:532:dfflibmap$9224;
    wire $auto$dfflibmap.cc:532:dfflibmap$9225;
    wire $auto$dfflibmap.cc:532:dfflibmap$9232;
    wire $auto$dfflibmap.cc:532:dfflibmap$9233;
    wire $auto$dfflibmap.cc:532:dfflibmap$9234;
    wire $auto$dfflibmap.cc:532:dfflibmap$9235;
    wire $auto$dfflibmap.cc:532:dfflibmap$9236;
    wire $auto$dfflibmap.cc:532:dfflibmap$9237;
    wire $auto$dfflibmap.cc:532:dfflibmap$9238;
    wire $auto$dfflibmap.cc:532:dfflibmap$9239;
    wire $auto$dfflibmap.cc:532:dfflibmap$9240;
    wire $auto$dfflibmap.cc:532:dfflibmap$9241;
    wire $auto$dfflibmap.cc:532:dfflibmap$9242;
    wire $auto$dfflibmap.cc:532:dfflibmap$9243;
    wire $auto$dfflibmap.cc:532:dfflibmap$9244;
    wire $auto$dfflibmap.cc:532:dfflibmap$9245;
    wire $auto$dfflibmap.cc:532:dfflibmap$9246;
    wire $auto$dfflibmap.cc:532:dfflibmap$9247;
    wire $auto$dfflibmap.cc:532:dfflibmap$9248;
    wire $auto$dfflibmap.cc:532:dfflibmap$9249;
    wire $auto$dfflibmap.cc:532:dfflibmap$9250;
    wire $auto$dfflibmap.cc:532:dfflibmap$9251;
    wire $auto$dfflibmap.cc:532:dfflibmap$9252;
    wire $auto$dfflibmap.cc:532:dfflibmap$9253;
    wire $auto$dfflibmap.cc:532:dfflibmap$9254;
    wire $auto$dfflibmap.cc:532:dfflibmap$9255;
    wire $auto$dfflibmap.cc:532:dfflibmap$9256;
    wire $auto$dfflibmap.cc:532:dfflibmap$9257;
    wire $auto$dfflibmap.cc:532:dfflibmap$9258;
    wire $auto$dfflibmap.cc:532:dfflibmap$9259;
    wire $auto$dfflibmap.cc:532:dfflibmap$9260;
    wire $auto$dfflibmap.cc:532:dfflibmap$9261;
    wire $auto$dfflibmap.cc:532:dfflibmap$9262;
    wire $auto$dfflibmap.cc:532:dfflibmap$9263;
    wire $auto$dfflibmap.cc:532:dfflibmap$9268;
    wire $auto$dfflibmap.cc:532:dfflibmap$9269;
    wire $auto$dfflibmap.cc:532:dfflibmap$9270;
    wire $auto$dfflibmap.cc:532:dfflibmap$9271;
    wire $auto$dfflibmap.cc:532:dfflibmap$9272;
    wire $auto$dfflibmap.cc:532:dfflibmap$9273;
    wire $auto$dfflibmap.cc:532:dfflibmap$9274;
    wire $auto$dfflibmap.cc:532:dfflibmap$9275;
    wire $auto$hilomap.cc:39:hilomap_worker$12030;
    wire [7:0] $flatten\CPU.$procmux$291.B;
    wire [215:0] $flatten\CPU.$procmux$415.B;
    wire [79:0] $flatten\CPU.$procmux$715.B;
    wire [7:0] CPU.ABH;
    wire [7:0] CPU.ABL;
    wire [7:0] CPU.ADD;
    wire CPU.ALU.AI7;
    wire CPU.ALU.BI7;
    wire CPU.ALU.CO;
    wire CPU.ALU.HC;
    wire CPU.ALU.N;
    wire [7:0] CPU.AXYS[0];
    wire [7:0] CPU.AXYS[1];
    wire [7:0] CPU.AXYS[2];
    wire [7:0] CPU.AXYS[3];
    wire CPU.C;
    wire CPU.D;
    wire [7:0] CPU.DIHOLD;
    wire [7:0] CPU.DIMUX;
    wire CPU.I;
    wire [7:0] CPU.IRHOLD;
    wire CPU.IRHOLD_valid;
    wire CPU.N;
    wire CPU.NMI_1;
    wire CPU.NMI_edge;
    wire [15:0] CPU.PC;
    wire CPU.V;
    wire CPU.Z;
    wire CPU.adc_bcd;
    wire CPU.adc_sbc;
    wire CPU.adj_bcd;
    wire CPU.backwards;
    wire CPU.bit_ins;
    wire CPU.clc;
    wire CPU.cld;
    wire CPU.cli;
    wire CPU.clv;
    wire CPU.compare;
    wire [2:0] CPU.cond_code;
    wire [1:0] CPU.dst_reg;
    wire CPU.inc;
    wire CPU.index_y;
    wire CPU.load_only;
    wire CPU.load_reg;
    wire [3:0] CPU.op;
    wire CPU.php;
    wire CPU.plp;
    wire CPU.res;
    wire CPU.rotate;
    wire CPU.sec;
    wire CPU.sed;
    wire CPU.sei;
    wire CPU.shift;
    wire CPU.shift_right;
    wire [1:0] CPU.src_reg;
    wire [5:0] CPU.state;
    wire CPU.store;
    wire CPU.write_back;
    wire cts_net_3116;
    wire cts_net_3117;
    wire cts_net_3118;
    wire cts_net_3119;
    wire cts_net_3120;
    wire cts_net_3121;
    wire cts_net_3122;
    wire cts_net_3123;
    wire cts_net_3124;
    wire cts_net_3125;
    wire cts_net_3126;
    wire cts_net_3127;
    wire cts_net_3128;
    wire cts_net_3129;
    wire cts_net_3130;
    wire cts_net_3131;
    wire cts_net_3132;
    wire cts_net_3133;
    wire cts_net_3134;
    wire cts_net_3135;
    wire cts_net_3136;
    wire cts_net_3137;
    wire cts_net_3138;
    wire cts_net_3139;
    wire cts_net_3140;
    wire cts_net_3141;
    wire cts_net_3142;
    wire cts_net_3143;
    wire cts_net_3144;
    wire cts_net_3145;
    wire cts_net_3146;
    wire cts_net_3147;
    wire cts_net_3148;
    wire cts_net_3149;
    wire cts_net_3150;
    wire cts_net_3151;
    wire cts_net_3152;
    wire cts_net_3153;
    wire cts_net_3154;
    wire cts_net_3155;
    wire cts_net_3156;
    wire cts_net_3157;
    wire cts_net_3158;
    wire cts_net_3159;
    wire cts_net_3160;
    wire cts_net_3161;
    wire cts_net_3162;
    wire cts_net_3163;
    wire cts_net_3164;
    wire cts_net_3165;
    wire cts_net_3166;
    wire cts_net_3167;
    wire cts_net_3168;
    wire cts_net_3169;
    wire cts_net_3170;
    wire cts_net_3171;
    wire cts_net_3172;
    wire cts_net_3173;
    wire cts_net_3174;
    wire cts_net_3175;
    wire cts_net_3176;
    wire cts_net_3177;
    wire cts_net_3178;
    wire cts_net_3179;
    wire cts_net_3180;
    wire cts_net_3181;
    wire cts_net_3182;
    wire cts_net_3183;
    wire cts_net_3184;
    wire cts_net_3185;
    wire cts_net_3186;
    wire cts_net_3187;
    wire cts_net_3188;
    wire cts_net_3189;
    wire cts_net_3190;
    wire cts_net_3191;
    wire cts_net_3192;
    wire cts_net_3193;
    wire cts_net_3194;
    wire cts_net_3195;
    wire cts_net_3196;
    wire cts_net_3197;
    wire cts_net_3198;
    wire cts_net_3199;
    wire cts_net_3200;
    wire cts_net_3201;
    wire cts_net_3202;
    wire cts_net_3203;

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10000 (
        .A($abc$9276$new_n1063), .B($abc$9276$new_n1068), .X($abc$9276$new_n1069)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10001 (
        .A($abc$9276$new_n1060), .B($abc$9276$new_n1069), .X($abc$9276$new_n1070)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10002 (
        .A($abc$9276$new_n1070), .Y($abc$9276$new_n1071)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10003 (
        .A($abc$9276$new_n1058), .B($abc$9276$new_n1071), .Y($abc$9276$new_n1072)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10004 (
        .A($abc$9276$new_n1051), .B($abc$9276$new_n1072), .Y($abc$9276$new_n1073)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10005 (
        .A($abc$9276$new_n1073), .Y($abc$9276$new_n1074)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10006 (
        .A($abc$9276$new_n1051), .B($abc$9276$new_n1072), .X($abc$9276$new_n1075)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10007 (
        .A($abc$9276$new_n1073), .B($abc$9276$new_n1075), .Y($abc$9276$new_n1076)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10008 (
        .A(in_35), .B($abc$9276$new_n1076), .Y($abc$9276$new_n1077)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10009 (
        .A(in_35), .B(CPU.PC), .X($abc$9276$new_n1078)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10010 (
        .A($abc$9276$new_n1077), .B($abc$9276$new_n1078), .Y($abc$9276$new_n1079)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10011 (
        .A($abc$9276$new_n1079), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8939)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10012 (
        .A(CPU.PC), .B($abc$9276$new_n1019), .Y($abc$9276$new_n1081)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10013 (
        .A(CPU.ADD), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1082)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10014 (
        .A(CPU.ADD), .B($abc$9276$new_n978), .Y($abc$9276$new_n1083)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10015 (
        .A($abc$9276$new_n1012), .B($abc$9276$new_n1083), .Y($abc$9276$new_n1084)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10016 (
        .A(CPU.ABL), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1085)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10017 (
        .A($abc$9276$new_n1082), .B($abc$9276$new_n1085), .Y($abc$9276$new_n1086)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10018 (
        .A($abc$9276$new_n1084), .B($abc$9276$new_n1086), .X($abc$9276$new_n1087)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10019 (
        .A($abc$9276$new_n1087), .Y($abc$9276$new_n1088)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10020 (
        .A($abc$9276$new_n1081), .B($abc$9276$new_n1088), .Y($abc$9276$new_n1089)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10021 (
        .A($abc$9276$new_n1074), .B($abc$9276$new_n1089), .Y($abc$9276$new_n1090)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10022 (
        .A($abc$9276$new_n1090), .Y($abc$9276$new_n1091)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10023 (
        .A($abc$9276$new_n1074), .B($abc$9276$new_n1089), .X($abc$9276$new_n1092)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10024 (
        .A($abc$9276$new_n1090), .B($abc$9276$new_n1092), .Y($abc$9276$new_n1093)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10025 (
        .A(in_35), .B($abc$9276$new_n1093), .Y($abc$9276$new_n1094)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10026 (
        .A(in_35), .B(CPU.PC), .X($abc$9276$new_n1095)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10027 (
        .A($abc$9276$new_n1094), .B($abc$9276$new_n1095), .Y($abc$9276$new_n1096)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10028 (
        .A($abc$9276$new_n1096), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8941)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10029 (
        .A(CPU.PC), .B($abc$9276$new_n1019), .Y($abc$9276$new_n1098)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10030 (
        .A(CPU.ADD), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1099)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10031 (
        .A($abc$9276$new_n375), .B($abc$9276$new_n977), .X($abc$9276$new_n1100)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10032 (
        .A($abc$9276$new_n1012), .B($abc$9276$new_n1100), .Y($abc$9276$new_n1101)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10033 (
        .A(CPU.ABL), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1102)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10034 (
        .A($abc$9276$new_n1099), .B($abc$9276$new_n1102), .Y($abc$9276$new_n1103)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10035 (
        .A($abc$9276$new_n1101), .B($abc$9276$new_n1103), .X($abc$9276$new_n1104)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10036 (
        .A($abc$9276$new_n1104), .Y($abc$9276$new_n1105)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10037 (
        .A($abc$9276$new_n1098), .B($abc$9276$new_n1105), .Y($abc$9276$new_n1106)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10038 (
        .A($abc$9276$new_n1091), .B($abc$9276$new_n1106), .Y($abc$9276$new_n1107)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10039 (
        .A($abc$9276$new_n1107), .Y($abc$9276$new_n1108)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10040 (
        .A($abc$9276$new_n1091), .B($abc$9276$new_n1106), .X($abc$9276$new_n1109)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10041 (
        .A($abc$9276$new_n1107), .B($abc$9276$new_n1109), .Y($abc$9276$new_n1110)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10042 (
        .A(in_35), .B($abc$9276$new_n1110), .Y($abc$9276$new_n1111)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10043 (
        .A(in_35), .B(CPU.PC), .X($abc$9276$new_n1112)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10044 (
        .A($abc$9276$new_n1111), .B($abc$9276$new_n1112), .Y($abc$9276$new_n1113)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10045 (
        .A($abc$9276$new_n1113), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8943)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10046 (
        .A(CPU.PC), .B($abc$9276$new_n1019), .Y($abc$9276$new_n1115)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10047 (
        .A(CPU.ADD), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1116)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10048 (
        .A(CPU.ADD), .B($abc$9276$new_n978), .Y($abc$9276$new_n1117)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10049 (
        .A(CPU.ABL), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1118)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10050 (
        .A($abc$9276$new_n1117), .B($abc$9276$new_n1118), .Y($abc$9276$new_n1119)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10051 (
        .A($abc$9276$new_n1119), .Y($abc$9276$new_n1120)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10052 (
        .A($abc$9276$new_n1116), .B($abc$9276$new_n1120), .Y($abc$9276$new_n1121)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10053 (
        .A($abc$9276$new_n1013), .B($abc$9276$new_n1121), .X($abc$9276$new_n1122)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10054 (
        .A($abc$9276$new_n1122), .Y($abc$9276$new_n1123)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10055 (
        .A($abc$9276$new_n1115), .B($abc$9276$new_n1123), .Y($abc$9276$new_n1124)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10056 (
        .A($abc$9276$new_n1108), .B($abc$9276$new_n1124), .Y($abc$9276$new_n1125)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10057 (
        .A($abc$9276$new_n1125), .Y($abc$9276$new_n1126)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10058 (
        .A($abc$9276$new_n1108), .B($abc$9276$new_n1124), .X($abc$9276$new_n1127)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10059 (
        .A($abc$9276$new_n1125), .B($abc$9276$new_n1127), .Y($abc$9276$new_n1128)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10060 (
        .A(in_35), .B(CPU.PC), .X($abc$9276$new_n1129)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10061 (
        .A(in_35), .B($abc$9276$new_n1128), .Y($abc$9276$new_n1130)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10062 (
        .A($abc$9276$new_n1129), .B($abc$9276$new_n1130), .Y($abc$9276$new_n1131)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10063 (
        .A($abc$9276$new_n1131), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8945)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10064 (
        .A(CPU.PC), .B($abc$9276$new_n1019), .Y($abc$9276$new_n1133)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10065 (
        .A(CPU.ADD), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1134)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10066 (
        .A($abc$9276$new_n376), .B($abc$9276$new_n977), .X($abc$9276$new_n1135)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10067 (
        .A($abc$9276$new_n1012), .B($abc$9276$new_n1135), .Y($abc$9276$new_n1136)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10068 (
        .A(CPU.ABL), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1137)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10069 (
        .A($abc$9276$new_n1134), .B($abc$9276$new_n1137), .Y($abc$9276$new_n1138)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10070 (
        .A($abc$9276$new_n1136), .B($abc$9276$new_n1138), .X($abc$9276$new_n1139)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10071 (
        .A($abc$9276$new_n1139), .Y($abc$9276$new_n1140)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10072 (
        .A($abc$9276$new_n1133), .B($abc$9276$new_n1140), .Y($abc$9276$new_n1141)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10073 (
        .A($abc$9276$new_n1126), .B($abc$9276$new_n1141), .Y($abc$9276$new_n1142)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10074 (
        .A($abc$9276$new_n1142), .Y($abc$9276$new_n1143)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10075 (
        .A($abc$9276$new_n1126), .B($abc$9276$new_n1141), .X($abc$9276$new_n1144)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10076 (
        .A($abc$9276$new_n1142), .B($abc$9276$new_n1144), .Y($abc$9276$new_n1145)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10077 (
        .A(in_35), .B($abc$9276$new_n1145), .Y($abc$9276$new_n1146)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10078 (
        .A(in_35), .B(CPU.PC), .X($abc$9276$new_n1147)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10079 (
        .A($abc$9276$new_n1146), .B($abc$9276$new_n1147), .Y($abc$9276$new_n1148)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10080 (
        .A($abc$9276$new_n1148), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8947)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10081 (
        .A(CPU.PC), .B($abc$9276$new_n1019), .Y($abc$9276$new_n1150)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10082 (
        .A(CPU.ALU.N), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1151)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10083 (
        .A($abc$9276$new_n372), .B($abc$9276$new_n977), .X($abc$9276$new_n1152)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10084 (
        .A($abc$9276$new_n1012), .B($abc$9276$new_n1152), .Y($abc$9276$new_n1153)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10085 (
        .A(CPU.ABL), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1154)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10086 (
        .A($abc$9276$new_n1151), .B($abc$9276$new_n1154), .Y($abc$9276$new_n1155)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10087 (
        .A($abc$9276$new_n1153), .B($abc$9276$new_n1155), .X($abc$9276$new_n1156)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10088 (
        .A($abc$9276$new_n1156), .Y($abc$9276$new_n1157)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10089 (
        .A($abc$9276$new_n1150), .B($abc$9276$new_n1157), .Y($abc$9276$new_n1158)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10090 (
        .A($abc$9276$new_n1143), .B($abc$9276$new_n1158), .Y($abc$9276$new_n1159)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10091 (
        .A($abc$9276$new_n1159), .Y($abc$9276$new_n1160)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10092 (
        .A($abc$9276$new_n1143), .B($abc$9276$new_n1158), .X($abc$9276$new_n1161)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10093 (
        .A($abc$9276$new_n1159), .B($abc$9276$new_n1161), .Y($abc$9276$new_n1162)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10094 (
        .A(in_35), .B(CPU.PC), .X($abc$9276$new_n1163)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10095 (
        .A(in_35), .B($abc$9276$new_n1162), .Y($abc$9276$new_n1164)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10096 (
        .A($abc$9276$new_n1163), .B($abc$9276$new_n1164), .Y($abc$9276$new_n1165)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10097 (
        .A($abc$9276$new_n1165), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8949)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10098 (
        .A(CPU.PC), .B($abc$9276$new_n1018), .Y($abc$9276$new_n1167)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10099 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1168)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10100 (
        .A(CPU.ABH), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1169)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10101 (
        .A(CPU.ABH), .B($abc$9276$new_n978), .Y($abc$9276$new_n1170)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10102 (
        .A($abc$9276$new_n1012), .B($abc$9276$new_n1170), .Y($abc$9276$new_n1171)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10103 (
        .A($abc$9276$new_n1171), .Y($abc$9276$new_n1172)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10104 (
        .A($abc$9276$new_n373), .B($abc$9276$new_n985), .X($abc$9276$new_n1173)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10105 (
        .A($abc$9276$new_n1169), .B($abc$9276$new_n1172), .Y($abc$9276$new_n1174)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10106 (
        .A($abc$9276$new_n1168), .B($abc$9276$new_n1173), .Y($abc$9276$new_n1175)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10107 (
        .A($abc$9276$new_n1174), .B($abc$9276$new_n1175), .X($abc$9276$new_n1176)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10108 (
        .A($abc$9276$new_n1176), .Y($abc$9276$new_n1177)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10109 (
        .A($abc$9276$new_n1167), .B($abc$9276$new_n1177), .Y($abc$9276$new_n1178)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10110 (
        .A($abc$9276$new_n1160), .B($abc$9276$new_n1178), .Y($abc$9276$new_n1179)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10111 (
        .A($abc$9276$new_n1179), .Y($abc$9276$new_n1180)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10112 (
        .A($abc$9276$new_n1160), .B($abc$9276$new_n1178), .X($abc$9276$new_n1181)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10113 (
        .A($abc$9276$new_n1179), .B($abc$9276$new_n1181), .Y($abc$9276$new_n1182)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10114 (
        .A(in_35), .B($abc$9276$new_n1182), .Y($abc$9276$new_n1183)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10115 (
        .A(in_35), .B(CPU.PC), .X($abc$9276$new_n1184)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10116 (
        .A($abc$9276$new_n1183), .B($abc$9276$new_n1184), .Y($abc$9276$new_n1185)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10117 (
        .A($abc$9276$new_n1185), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8951)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10118 (
        .A(CPU.PC), .B($abc$9276$new_n1018), .Y($abc$9276$new_n1187)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10119 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1188)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10120 (
        .A(CPU.ABH), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1189)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10121 (
        .A(CPU.ABH), .B($abc$9276$new_n978), .Y($abc$9276$new_n1190)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10122 (
        .A(CPU.ADD), .B($abc$9276$new_n986), .Y($abc$9276$new_n1191)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10123 (
        .A($abc$9276$new_n1189), .B($abc$9276$new_n1190), .Y($abc$9276$new_n1192)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10124 (
        .A($abc$9276$new_n1013), .B($abc$9276$new_n1192), .X($abc$9276$new_n1193)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10125 (
        .A($abc$9276$new_n1188), .B($abc$9276$new_n1191), .Y($abc$9276$new_n1194)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10126 (
        .A($abc$9276$new_n1193), .B($abc$9276$new_n1194), .X($abc$9276$new_n1195)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10127 (
        .A($abc$9276$new_n1195), .Y($abc$9276$new_n1196)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10128 (
        .A($abc$9276$new_n1187), .B($abc$9276$new_n1196), .Y($abc$9276$new_n1197)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10129 (
        .A($abc$9276$new_n1180), .B($abc$9276$new_n1197), .Y($abc$9276$new_n1198)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10130 (
        .A($abc$9276$new_n1198), .Y($abc$9276$new_n1199)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10131 (
        .A($abc$9276$new_n1180), .B($abc$9276$new_n1197), .X($abc$9276$new_n1200)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10132 (
        .A($abc$9276$new_n1198), .B($abc$9276$new_n1200), .Y($abc$9276$new_n1201)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10133 (
        .A(in_35), .B($abc$9276$new_n1201), .Y($abc$9276$new_n1202)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10134 (
        .A(in_35), .B(CPU.PC), .X($abc$9276$new_n1203)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10135 (
        .A($abc$9276$new_n1202), .B($abc$9276$new_n1203), .Y($abc$9276$new_n1204)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10136 (
        .A($abc$9276$new_n1204), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8953)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10137 (
        .A(CPU.PC), .B($abc$9276$new_n1018), .Y($abc$9276$new_n1206)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10138 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1207)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10139 (
        .A(CPU.ABH), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1208)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10140 (
        .A($abc$9276$new_n374), .B($abc$9276$new_n985), .X($abc$9276$new_n1209)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10141 (
        .A(CPU.ABH), .B($abc$9276$new_n978), .Y($abc$9276$new_n1210)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10142 (
        .A($abc$9276$new_n1210), .Y($abc$9276$new_n1211)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10143 (
        .A($abc$9276$new_n1012), .B($abc$9276$new_n1208), .Y($abc$9276$new_n1212)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10144 (
        .A($abc$9276$new_n1211), .B($abc$9276$new_n1212), .X($abc$9276$new_n1213)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10145 (
        .A($abc$9276$new_n1207), .B($abc$9276$new_n1209), .Y($abc$9276$new_n1214)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10146 (
        .A($abc$9276$new_n1213), .B($abc$9276$new_n1214), .X($abc$9276$new_n1215)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10147 (
        .A($abc$9276$new_n1215), .Y($abc$9276$new_n1216)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10148 (
        .A($abc$9276$new_n1206), .B($abc$9276$new_n1216), .Y($abc$9276$new_n1217)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10149 (
        .A($abc$9276$new_n1199), .B($abc$9276$new_n1217), .Y($abc$9276$new_n1218)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10150 (
        .A($abc$9276$new_n1218), .Y($abc$9276$new_n1219)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10151 (
        .A($abc$9276$new_n1199), .B($abc$9276$new_n1217), .X($abc$9276$new_n1220)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10152 (
        .A($abc$9276$new_n1218), .B($abc$9276$new_n1220), .Y($abc$9276$new_n1221)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10153 (
        .A(in_35), .B(CPU.PC), .X($abc$9276$new_n1222)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10154 (
        .A(in_35), .B($abc$9276$new_n1221), .Y($abc$9276$new_n1223)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10155 (
        .A($abc$9276$new_n1222), .B($abc$9276$new_n1223), .Y($abc$9276$new_n1224)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10156 (
        .A($abc$9276$new_n1224), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8955)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10157 (
        .A(CPU.PC), .B($abc$9276$new_n1018), .Y($abc$9276$new_n1226)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10158 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1227)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10159 (
        .A(CPU.ABH), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1228)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10160 (
        .A(CPU.ADD), .B($abc$9276$new_n986), .Y($abc$9276$new_n1229)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10161 (
        .A(CPU.ABH), .B($abc$9276$new_n978), .Y($abc$9276$new_n1230)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10162 (
        .A($abc$9276$new_n1229), .B($abc$9276$new_n1230), .Y($abc$9276$new_n1231)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10163 (
        .A($abc$9276$new_n1013), .B($abc$9276$new_n1231), .X($abc$9276$new_n1232)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10164 (
        .A($abc$9276$new_n1227), .B($abc$9276$new_n1228), .Y($abc$9276$new_n1233)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10165 (
        .A($abc$9276$new_n1232), .B($abc$9276$new_n1233), .X($abc$9276$new_n1234)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10166 (
        .A($abc$9276$new_n1234), .Y($abc$9276$new_n1235)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10167 (
        .A($abc$9276$new_n1226), .B($abc$9276$new_n1235), .Y($abc$9276$new_n1236)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10168 (
        .A($abc$9276$new_n1219), .B($abc$9276$new_n1236), .Y($abc$9276$new_n1237)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10169 (
        .A($abc$9276$new_n1237), .Y($abc$9276$new_n1238)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10170 (
        .A($abc$9276$new_n1219), .B($abc$9276$new_n1236), .X($abc$9276$new_n1239)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10171 (
        .A($abc$9276$new_n1237), .B($abc$9276$new_n1239), .Y($abc$9276$new_n1240)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10172 (
        .A(in_35), .B($abc$9276$new_n1240), .Y($abc$9276$new_n1241)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10173 (
        .A(in_35), .B(CPU.PC), .X($abc$9276$new_n1242)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10174 (
        .A($abc$9276$new_n1241), .B($abc$9276$new_n1242), .Y($abc$9276$new_n1243)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10175 (
        .A($abc$9276$new_n1243), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8957)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10176 (
        .A(CPU.PC), .B($abc$9276$new_n1018), .Y($abc$9276$new_n1245)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10177 (
        .A($abc$9276$new_n1245), .Y($abc$9276$new_n1246)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10178 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1247)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10179 (
        .A($abc$9276$new_n1247), .Y($abc$9276$new_n1248)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10180 (
        .A(CPU.ABH), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1249)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10181 (
        .A($abc$9276$new_n375), .B($abc$9276$new_n985), .X($abc$9276$new_n1250)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10182 (
        .A(CPU.ABH), .B($abc$9276$new_n978), .Y($abc$9276$new_n1251)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10183 (
        .A($abc$9276$new_n1251), .Y($abc$9276$new_n1252)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10184 (
        .A($abc$9276$new_n1249), .B($abc$9276$new_n1250), .Y($abc$9276$new_n1253)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10185 (
        .A($abc$9276$new_n1252), .B($abc$9276$new_n1253), .X($abc$9276$new_n1254)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10186 (
        .A($abc$9276$new_n1248), .B($abc$9276$new_n1254), .X($abc$9276$new_n1255)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10187 (
        .A($abc$9276$new_n1013), .B($abc$9276$new_n1255), .X($abc$9276$new_n1256)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10188 (
        .A($abc$9276$new_n1246), .B($abc$9276$new_n1256), .X($abc$9276$new_n1257)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10189 (
        .A($abc$9276$new_n1238), .B($abc$9276$new_n1257), .Y($abc$9276$new_n1258)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10190 (
        .A($abc$9276$new_n1258), .Y($abc$9276$new_n1259)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10191 (
        .A($abc$9276$new_n1238), .B($abc$9276$new_n1257), .X($abc$9276$new_n1260)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10192 (
        .A($abc$9276$new_n1258), .B($abc$9276$new_n1260), .Y($abc$9276$new_n1261)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10193 (
        .A(in_35), .B($abc$9276$new_n1261), .Y($abc$9276$new_n1262)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10194 (
        .A(in_35), .B(CPU.PC), .X($abc$9276$new_n1263)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10195 (
        .A($abc$9276$new_n1262), .B($abc$9276$new_n1263), .Y($abc$9276$new_n1264)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10196 (
        .A($abc$9276$new_n1264), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8959)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10197 (
        .A(CPU.PC), .B($abc$9276$new_n1018), .Y($abc$9276$new_n1266)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10198 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1267)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10199 (
        .A($abc$9276$new_n1267), .Y($abc$9276$new_n1268)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10200 (
        .A(CPU.ABH), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1269)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10201 (
        .A(CPU.ABH), .B($abc$9276$new_n978), .Y($abc$9276$new_n1270)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10202 (
        .A($abc$9276$new_n1012), .B($abc$9276$new_n1270), .Y($abc$9276$new_n1271)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10203 (
        .A(CPU.ADD), .B($abc$9276$new_n986), .Y($abc$9276$new_n1272)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10204 (
        .A($abc$9276$new_n1269), .B($abc$9276$new_n1272), .Y($abc$9276$new_n1273)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10205 (
        .A($abc$9276$new_n1271), .B($abc$9276$new_n1273), .X($abc$9276$new_n1274)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10206 (
        .A($abc$9276$new_n1274), .Y($abc$9276$new_n1275)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10207 (
        .A($abc$9276$new_n1266), .B($abc$9276$new_n1275), .Y($abc$9276$new_n1276)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10208 (
        .A($abc$9276$new_n1268), .B($abc$9276$new_n1276), .X($abc$9276$new_n1277)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10209 (
        .A($abc$9276$new_n1259), .B($abc$9276$new_n1277), .Y($abc$9276$new_n1278)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10210 (
        .A($abc$9276$new_n1278), .Y($abc$9276$new_n1279)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10211 (
        .A($abc$9276$new_n1259), .B($abc$9276$new_n1277), .X($abc$9276$new_n1280)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10212 (
        .A($abc$9276$new_n1278), .B($abc$9276$new_n1280), .Y($abc$9276$new_n1281)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10213 (
        .A(in_35), .B($abc$9276$new_n1281), .Y($abc$9276$new_n1282)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10214 (
        .A(in_35), .B(CPU.PC), .X($abc$9276$new_n1283)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10215 (
        .A($abc$9276$new_n1282), .B($abc$9276$new_n1283), .Y($abc$9276$new_n1284)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10216 (
        .A($abc$9276$new_n1284), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8961)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10217 (
        .A(CPU.PC), .B($abc$9276$new_n1018), .Y($abc$9276$new_n1286)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10218 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1287)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10219 (
        .A(CPU.ABH), .B($abc$9276$new_n978), .Y($abc$9276$new_n1288)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10220 (
        .A($abc$9276$new_n376), .B($abc$9276$new_n985), .X($abc$9276$new_n1289)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10221 (
        .A($abc$9276$new_n1288), .B($abc$9276$new_n1289), .Y($abc$9276$new_n1290)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10222 (
        .A($abc$9276$new_n1013), .B($abc$9276$new_n1290), .X($abc$9276$new_n1291)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10223 (
        .A(CPU.ABH), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1292)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10224 (
        .A($abc$9276$new_n1287), .B($abc$9276$new_n1292), .Y($abc$9276$new_n1293)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10225 (
        .A($abc$9276$new_n1291), .B($abc$9276$new_n1293), .X($abc$9276$new_n1294)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10226 (
        .A($abc$9276$new_n1294), .Y($abc$9276$new_n1295)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10227 (
        .A($abc$9276$new_n1286), .B($abc$9276$new_n1295), .Y($abc$9276$new_n1296)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10228 (
        .A($abc$9276$new_n1279), .B($abc$9276$new_n1296), .Y($abc$9276$new_n1297)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10229 (
        .A($abc$9276$new_n1279), .B($abc$9276$new_n1296), .X($abc$9276$new_n1298)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10230 (
        .A($abc$9276$new_n1297), .B($abc$9276$new_n1298), .Y($abc$9276$new_n1299)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10231 (
        .A(in_35), .B($abc$9276$new_n1299), .Y($abc$9276$new_n1300)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10232 (
        .A(in_35), .B(CPU.PC), .X($abc$9276$new_n1301)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10233 (
        .A($abc$9276$new_n1300), .B($abc$9276$new_n1301), .Y($abc$9276$new_n1302)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10234 (
        .A($abc$9276$new_n1302), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8963)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10235 (
        .A(CPU.PC), .B($abc$9276$new_n1018), .Y($abc$9276$new_n1304)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10236 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1305)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10237 (
        .A(CPU.ABH), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1306)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10238 (
        .A($abc$9276$new_n372), .B($abc$9276$new_n985), .X($abc$9276$new_n1307)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10239 (
        .A(CPU.ABH), .B($abc$9276$new_n978), .Y($abc$9276$new_n1308)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10240 (
        .A($abc$9276$new_n1305), .B($abc$9276$new_n1307), .Y($abc$9276$new_n1309)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10241 (
        .A($abc$9276$new_n1306), .B($abc$9276$new_n1308), .Y($abc$9276$new_n1310)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10242 (
        .A($abc$9276$new_n1013), .B($abc$9276$new_n1310), .X($abc$9276$new_n1311)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10243 (
        .A($abc$9276$new_n1309), .B($abc$9276$new_n1311), .X($abc$9276$new_n1312)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10244 (
        .A($abc$9276$new_n1312), .Y($abc$9276$new_n1313)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10245 (
        .A($abc$9276$new_n1304), .B($abc$9276$new_n1313), .Y($abc$9276$new_n1314)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10246 (
        .A($abc$9276$new_n1297), .B($abc$9276$new_n1314), .X($abc$9276$new_n1315)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10247 (
        .A($abc$9276$new_n1297), .B($abc$9276$new_n1314), .Y($abc$9276$new_n1316)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10248 (
        .A($abc$9276$new_n359), .B(CPU.PC), .Y($abc$9276$new_n1317)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10249 (
        .A($abc$9276$new_n1315), .B($abc$9276$new_n1316), .Y($abc$9276$new_n1318)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10250 (
        .A(in_35), .B($abc$9276$new_n1318), .Y($abc$9276$new_n1319)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10251 (
        .A($abc$9276$new_n1317), .B($abc$9276$new_n1319), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8965)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10252 (
        .A($abc$9276$new_n359), .B(CPU.cond_code), .Y($abc$9276$new_n1321)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10253 (
        .A(in_35), .B($abc$9276$new_n827), .Y($abc$9276$new_n1322)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10254 (
        .A($abc$9276$new_n1321), .B($abc$9276$new_n1322), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8971)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10255 (
        .A($abc$9276$new_n359), .B(CPU.cond_code), .Y($abc$9276$new_n1324)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10256 (
        .A(in_35), .B($abc$9276$new_n789), .Y($abc$9276$new_n1325)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10257 (
        .A($abc$9276$new_n1324), .B($abc$9276$new_n1325), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8973)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10258 (
        .A($abc$9276$new_n359), .B(CPU.cond_code), .Y($abc$9276$new_n1327)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10259 (
        .A(in_35), .B($abc$9276$new_n779), .Y($abc$9276$new_n1328)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10260 (
        .A($abc$9276$new_n1327), .B($abc$9276$new_n1328), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8975)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10261 (
        .A(CPU.cld), .B(CPU.sed), .X($abc$9276$new_n1330)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10262 (
        .A(CPU.cld), .B($abc$9276$new_n377), .Y($abc$9276$new_n1331)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10263 (
        .A(oeb_16), .B(CPU.sed), .Y($abc$9276$new_n1332)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10264 (
        .A($abc$9276$new_n354), .B($abc$9276$new_n1332), .Y($abc$9276$new_n1333)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10265 (
        .A($abc$9276$new_n1331), .B($abc$9276$new_n1333), .Y($abc$9276$new_n1334)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10266 (
        .A(CPU.plp), .B($abc$9276$new_n1334), .X($abc$9276$new_n1335)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10267 (
        .A(CPU.plp), .B(CPU.ADD), .Y($abc$9276$new_n1336)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10268 (
        .A($abc$9276$new_n1335), .B($abc$9276$new_n1336), .Y($abc$9276$new_n1337)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10269 (
        .A($abc$9276$new_n732), .B($abc$9276$new_n1337), .Y($abc$9276$new_n1338)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10270 (
        .A($abc$9276$new_n545), .B($abc$9276$new_n729), .X($abc$9276$new_n1339)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10271 (
        .A($abc$9276$new_n1339), .Y($abc$9276$new_n1340)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10272 (
        .A($abc$9276$new_n429), .B($abc$9276$new_n1330), .Y($abc$9276$new_n1341)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10273 (
        .A(CPU.D), .B($abc$9276$new_n729), .Y($abc$9276$new_n1342)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10274 (
        .A($abc$9276$new_n742), .B($abc$9276$new_n1341), .Y($abc$9276$new_n1343)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10275 (
        .A($abc$9276$new_n1342), .B($abc$9276$new_n1343), .X($abc$9276$new_n1344)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10276 (
        .A($abc$9276$new_n1338), .B($abc$9276$new_n1344), .Y($abc$9276$new_n1345)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10277 (
        .A($abc$9276$new_n1340), .B($abc$9276$new_n1345), .X($abc$9276$auto$rtlil.cc:3205:MuxGate$8981)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10278 (
        .A(CPU.load_reg), .B($abc$9276$new_n658), .Y($abc$9276$new_n1347)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10279 (
        .A($abc$9276$new_n358), .B($abc$9276$new_n1347), .Y($abc$9276$new_n1348)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10280 (
        .A($abc$9276$new_n429), .B($abc$9276$new_n1348), .Y($abc$9276$new_n1349)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10281 (
        .A($abc$9276$new_n742), .B($abc$9276$new_n1349), .Y($abc$9276$new_n1350)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10282 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n420), .X($abc$9276$new_n1351)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10283 (
        .A($abc$9276$new_n1351), .Y($abc$9276$new_n1352)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10284 (
        .A($abc$9276$new_n729), .B($abc$9276$new_n1351), .Y($abc$9276$new_n1353)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10285 (
        .A($abc$9276$new_n1353), .Y($abc$9276$new_n1354)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10286 (
        .A($abc$9276$new_n739), .B($abc$9276$new_n1354), .Y($abc$9276$new_n1355)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10287 (
        .A($abc$9276$new_n361), .B($abc$9276$new_n1355), .X($abc$9276$new_n1356)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10288 (
        .A($abc$9276$new_n1350), .B($abc$9276$new_n1356), .X($abc$9276$new_n1357)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10289 (
        .A($abc$9276$new_n372), .B($abc$9276$new_n1351), .X($abc$9276$new_n1358)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10290 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1351), .Y($abc$9276$new_n1359)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10291 (
        .A($abc$9276$new_n741), .B($abc$9276$new_n1359), .X($abc$9276$new_n1360)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10292 (
        .A($abc$9276$new_n1358), .B($abc$9276$new_n1360), .Y($abc$9276$new_n1361)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10293 (
        .A(CPU.ALU.N), .B($abc$9276$new_n1350), .Y($abc$9276$new_n1362)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10294 (
        .A($abc$9276$new_n1353), .B($abc$9276$new_n1362), .X($abc$9276$new_n1363)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10295 (
        .A($abc$9276$new_n1357), .B($abc$9276$new_n1363), .Y($abc$9276$new_n1364)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10296 (
        .A($abc$9276$new_n1361), .B($abc$9276$new_n1364), .X($abc$9276$auto$rtlil.cc:3205:MuxGate$8983)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10297 (
        .A($abc$9276$new_n505), .B($abc$9276$new_n729), .X($abc$9276$new_n1366)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10298 (
        .A(CPU.plp), .B(CPU.ADD), .Y($abc$9276$new_n1367)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10299 (
        .A(CPU.bit_ins), .B($abc$9276$new_n1348), .X($abc$9276$new_n1368)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10300 (
        .A(CPU.ADD), .B(CPU.ADD), .X($abc$9276$new_n1369)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10301 (
        .A(CPU.ADD), .B(CPU.ADD), .X($abc$9276$new_n1370)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10302 (
        .A($abc$9276$new_n1369), .B($abc$9276$new_n1370), .X($abc$9276$new_n1371)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10303 (
        .A(CPU.ALU.N), .B(CPU.ADD), .X($abc$9276$new_n1372)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10304 (
        .A(CPU.ADD), .B(CPU.ADD), .X($abc$9276$new_n1373)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10305 (
        .A($abc$9276$new_n1372), .B($abc$9276$new_n1373), .X($abc$9276$new_n1374)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10306 (
        .A($abc$9276$new_n1371), .B($abc$9276$new_n1374), .X($abc$9276$new_n1375)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10307 (
        .A(CPU.plp), .B($abc$9276$new_n1375), .X($abc$9276$new_n1376)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10308 (
        .A($abc$9276$new_n1376), .Y($abc$9276$new_n1377)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10309 (
        .A($abc$9276$new_n1368), .B($abc$9276$new_n1377), .Y($abc$9276$new_n1378)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10310 (
        .A($abc$9276$new_n1367), .B($abc$9276$new_n1378), .Y($abc$9276$new_n1379)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10311 (
        .A($abc$9276$new_n732), .B($abc$9276$new_n1379), .Y($abc$9276$new_n1380)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10312 (
        .A($abc$9276$new_n1366), .B($abc$9276$new_n1380), .Y($abc$9276$new_n1381)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10313 (
        .A($abc$9276$new_n1351), .B($abc$9276$new_n1381), .Y($abc$9276$new_n1382)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10314 (
        .A($abc$9276$new_n1351), .B($abc$9276$new_n1375), .X($abc$9276$new_n1383)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10315 (
        .A($abc$9276$new_n429), .B($abc$9276$new_n1368), .Y($abc$9276$new_n1384)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10316 (
        .A(CPU.Z), .B($abc$9276$new_n742), .Y($abc$9276$new_n1385)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10317 (
        .A($abc$9276$new_n1353), .B($abc$9276$new_n1385), .X($abc$9276$new_n1386)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10318 (
        .A($abc$9276$new_n1386), .Y($abc$9276$new_n1387)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10319 (
        .A($abc$9276$new_n1384), .B($abc$9276$new_n1387), .Y($abc$9276$new_n1388)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10320 (
        .A($abc$9276$new_n1383), .B($abc$9276$new_n1388), .Y($abc$9276$new_n1389)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10321 (
        .A($abc$9276$new_n1389), .Y($abc$9276$new_n1390)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10322 (
        .A($abc$9276$new_n1382), .B($abc$9276$new_n1390), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8989)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10323 (
        .A(CPU.shift), .B($abc$9276$new_n1352), .Y($abc$9276$new_n1392)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10324 (
        .A($abc$9276$new_n1392), .Y($abc$9276$new_n1393)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10325 (
        .A($abc$9276$new_n730), .B($abc$9276$new_n1392), .Y($abc$9276$new_n1394)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10326 (
        .A(CPU.compare), .B(CPU.shift), .X($abc$9276$new_n1395)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10327 (
        .A(CPU.adc_sbc), .B($abc$9276$new_n1395), .X($abc$9276$new_n1396)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10328 (
        .A($abc$9276$new_n1396), .Y($abc$9276$new_n1397)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10329 (
        .A($abc$9276$new_n1394), .B($abc$9276$new_n1396), .Y($abc$9276$new_n1398)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10330 (
        .A(CPU.ALU.CO), .B($abc$9276$new_n1398), .X($abc$9276$new_n1399)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10331 (
        .A(oeb_16), .B(CPU.sec), .Y($abc$9276$new_n1400)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10332 (
        .A(CPU.clc), .B(oeb_0), .Y($abc$9276$new_n1401)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10333 (
        .A(CPU.clc), .B($abc$9276$new_n1400), .X($abc$9276$new_n1402)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10334 (
        .A($abc$9276$new_n1401), .B($abc$9276$new_n1402), .Y($abc$9276$new_n1403)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10335 (
        .A(CPU.plp), .B($abc$9276$new_n1403), .X($abc$9276$new_n1404)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10336 (
        .A(CPU.plp), .B($abc$9276$new_n373), .Y($abc$9276$new_n1405)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10337 (
        .A($abc$9276$new_n1404), .B($abc$9276$new_n1405), .Y($abc$9276$new_n1406)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10338 (
        .A($abc$9276$new_n1397), .B($abc$9276$new_n1406), .Y($abc$9276$new_n1407)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10339 (
        .A($flatten\CPU.$procmux$415.B), .B($abc$9276$new_n429), .Y($abc$9276$new_n1408)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10340 (
        .A($abc$9276$new_n1408), .Y($abc$9276$new_n1409)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10341 (
        .A($abc$9276$new_n1407), .B($abc$9276$new_n1409), .Y($abc$9276$new_n1410)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10342 (
        .A($abc$9276$new_n730), .B($abc$9276$new_n1410), .X($abc$9276$new_n1411)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10343 (
        .A($abc$9276$new_n487), .B($abc$9276$new_n729), .X($abc$9276$new_n1412)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10344 (
        .A($abc$9276$new_n1392), .B($abc$9276$new_n1412), .Y($abc$9276$new_n1413)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10345 (
        .A($abc$9276$new_n1413), .Y($abc$9276$new_n1414)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10346 (
        .A($abc$9276$new_n1411), .B($abc$9276$new_n1414), .Y($abc$9276$new_n1415)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10347 (
        .A($abc$9276$new_n1399), .B($abc$9276$new_n1415), .Y($abc$9276$new_n1416)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10348 (
        .A(CPU.plp), .B(CPU.clc), .X($abc$9276$new_n1417)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10349 (
        .A(CPU.sec), .B($abc$9276$new_n1417), .X($abc$9276$new_n1418)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10350 (
        .A($abc$9276$new_n1396), .B($abc$9276$new_n1418), .X($abc$9276$new_n1419)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10351 (
        .A($abc$9276$new_n1409), .B($abc$9276$new_n1419), .Y($abc$9276$new_n1420)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10352 (
        .A(CPU.C), .B($abc$9276$new_n729), .Y($abc$9276$new_n1421)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10353 (
        .A($abc$9276$new_n1421), .Y($abc$9276$new_n1422)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10354 (
        .A($abc$9276$new_n1420), .B($abc$9276$new_n1422), .Y($abc$9276$new_n1423)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10355 (
        .A($abc$9276$new_n1393), .B($abc$9276$new_n1423), .X($abc$9276$new_n1424)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10356 (
        .A($abc$9276$new_n1416), .B($abc$9276$new_n1424), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8991)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10357 (
        .A($abc$9276$new_n359), .B(CPU.backwards), .Y($abc$9276$new_n1426)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10358 (
        .A($abc$9276$new_n624), .B($abc$9276$new_n1426), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8993)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10359 (
        .A($abc$9276$new_n348), .B($abc$9276$new_n449), .X($abc$9276$new_n1428)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10360 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n449), .Y($abc$9276$new_n1429)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10361 (
        .A($abc$9276$new_n1428), .B($abc$9276$new_n1429), .Y($abc$9276$new_n1430)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10362 (
        .A($abc$9276$new_n467), .B($abc$9276$new_n1430), .Y($abc$9276$new_n1431)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10363 (
        .A($abc$9276$new_n347), .B($abc$9276$new_n449), .X($abc$9276$new_n1432)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10364 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n449), .Y($abc$9276$new_n1433)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10365 (
        .A($abc$9276$new_n1432), .B($abc$9276$new_n1433), .Y($abc$9276$new_n1434)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10366 (
        .A($abc$9276$new_n466), .B($abc$9276$new_n1434), .Y($abc$9276$new_n1435)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10367 (
        .A($abc$9276$new_n1431), .B($abc$9276$new_n1435), .Y($abc$9276$new_n1436)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10368 (
        .A($abc$9276$new_n406), .B($abc$9276$new_n1436), .Y($abc$9276$new_n1437)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10369 (
        .A($abc$9276$new_n393), .B($abc$9276$new_n415), .X($abc$9276$new_n1438)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10370 (
        .A($abc$9276$new_n383), .B($abc$9276$new_n399), .X($abc$9276$new_n1439)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10371 (
        .A($abc$9276$new_n432), .B($abc$9276$new_n1439), .X($abc$9276$new_n1440)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10372 (
        .A($abc$9276$new_n1438), .B($abc$9276$new_n1440), .Y($abc$9276$new_n1441)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10373 (
        .A($abc$9276$new_n388), .B($abc$9276$new_n431), .X($abc$9276$new_n1442)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10374 (
        .A($abc$9276$new_n435), .B($abc$9276$new_n1442), .Y($abc$9276$new_n1443)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10375 (
        .A($abc$9276$new_n1441), .B($abc$9276$new_n1443), .X($abc$9276$new_n1444)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10376 (
        .A($abc$9276$new_n729), .B($abc$9276$new_n1012), .Y($abc$9276$new_n1445)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10377 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n976), .X($abc$9276$new_n1446)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10378 (
        .A($abc$9276$new_n388), .B($abc$9276$new_n409), .X($abc$9276$new_n1447)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10379 (
        .A($abc$9276$new_n1446), .B($abc$9276$new_n1447), .Y($abc$9276$new_n1448)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10380 (
        .A($abc$9276$new_n1445), .B($abc$9276$new_n1448), .X($abc$9276$new_n1449)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10381 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n409), .X($abc$9276$new_n1450)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10382 (
        .A($abc$9276$new_n1450), .Y($abc$9276$new_n1451)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10383 (
        .A($abc$9276$new_n413), .B($abc$9276$new_n1450), .Y($abc$9276$new_n1452)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10384 (
        .A($abc$9276$new_n393), .B($abc$9276$new_n995), .X($abc$9276$new_n1453)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10385 (
        .A($abc$9276$new_n1453), .Y($abc$9276$new_n1454)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10386 (
        .A($abc$9276$new_n419), .B($abc$9276$new_n1452), .X($abc$9276$new_n1455)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10387 (
        .A($abc$9276$new_n1449), .B($abc$9276$new_n1454), .X($abc$9276$new_n1456)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10388 (
        .A($abc$9276$new_n1455), .B($abc$9276$new_n1456), .X($abc$9276$new_n1457)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10389 (
        .A($abc$9276$new_n1457), .Y($abc$9276$new_n1458)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10390 (
        .A($abc$9276$new_n393), .B($abc$9276$new_n434), .X($abc$9276$new_n1459)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10391 (
        .A($abc$9276$new_n395), .B($abc$9276$new_n400), .X($abc$9276$new_n1460)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10392 (
        .A($abc$9276$new_n388), .B($abc$9276$new_n1460), .X($abc$9276$new_n1461)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10393 (
        .A($abc$9276$new_n1459), .B($abc$9276$new_n1461), .Y($abc$9276$new_n1462)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10394 (
        .A($abc$9276$new_n388), .B($abc$9276$new_n1439), .X($abc$9276$new_n1463)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10395 (
        .A($abc$9276$new_n393), .B($abc$9276$new_n1439), .X($abc$9276$new_n1464)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10396 (
        .A($abc$9276$new_n1463), .B($abc$9276$new_n1464), .Y($abc$9276$new_n1465)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10397 (
        .A($abc$9276$new_n1462), .B($abc$9276$new_n1465), .X($abc$9276$new_n1466)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10398 (
        .A($abc$9276$new_n1000), .B($abc$9276$new_n1466), .X($abc$9276$new_n1467)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10399 (
        .A($abc$9276$new_n1444), .B($abc$9276$new_n1467), .X($abc$9276$new_n1468)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10400 (
        .A($abc$9276$new_n1457), .B($abc$9276$new_n1468), .X($abc$9276$new_n1469)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10401 (
        .A($abc$9276$new_n388), .B($abc$9276$new_n401), .X($abc$9276$new_n1470)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10402 (
        .A($abc$9276$new_n1470), .Y($abc$9276$new_n1471)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10403 (
        .A($abc$9276$new_n393), .B($abc$9276$new_n1460), .X($abc$9276$new_n1472)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10404 (
        .A($abc$9276$new_n985), .B($abc$9276$new_n1472), .Y($abc$9276$new_n1473)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10405 (
        .A($abc$9276$new_n1471), .B($abc$9276$new_n1473), .X($abc$9276$new_n1474)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10406 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n1460), .X($abc$9276$new_n1475)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10407 (
        .A($abc$9276$new_n1475), .Y($abc$9276$new_n1476)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10408 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n434), .X($abc$9276$new_n1477)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10409 (
        .A($abc$9276$new_n1475), .B($abc$9276$new_n1477), .Y($abc$9276$new_n1478)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10410 (
        .A($abc$9276$new_n1352), .B($abc$9276$new_n1478), .X($abc$9276$new_n1479)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10411 (
        .A($abc$9276$new_n1474), .B($abc$9276$new_n1479), .X($abc$9276$new_n1480)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10412 (
        .A($abc$9276$new_n384), .B($abc$9276$new_n388), .X($abc$9276$new_n1481)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10413 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n415), .X($abc$9276$new_n1482)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10414 (
        .A($abc$9276$new_n1481), .B($abc$9276$new_n1482), .Y($abc$9276$new_n1483)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10415 (
        .A($abc$9276$new_n978), .B($abc$9276$new_n1483), .X($abc$9276$new_n1484)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10416 (
        .A($abc$9276$new_n406), .B($abc$9276$new_n1484), .X($abc$9276$new_n1485)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10417 (
        .A($abc$9276$new_n1480), .B($abc$9276$new_n1485), .X($abc$9276$new_n1486)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10418 (
        .A($abc$9276$new_n1469), .B($abc$9276$new_n1486), .X($abc$9276$new_n1487)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10419 (
        .A($abc$9276$new_n1487), .Y($abc$9276$new_n1488)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10420 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1489)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10421 (
        .A(CPU.ADD), .B($abc$9276$new_n1469), .Y($abc$9276$new_n1490)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10422 (
        .A(CPU.ABL), .B($abc$9276$new_n1480), .Y($abc$9276$new_n1491)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10423 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1483), .Y($abc$9276$new_n1492)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10424 (
        .A($abc$9276$new_n1025), .B($abc$9276$new_n1492), .Y($abc$9276$new_n1493)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10425 (
        .A($abc$9276$new_n1493), .Y($abc$9276$new_n1494)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10426 (
        .A($abc$9276$new_n1491), .B($abc$9276$new_n1494), .Y($abc$9276$new_n1495)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10427 (
        .A($abc$9276$new_n1495), .Y($abc$9276$new_n1496)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10428 (
        .A($abc$9276$new_n1490), .B($abc$9276$new_n1496), .Y($abc$9276$new_n1497)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10429 (
        .A($abc$9276$new_n1497), .Y($abc$9276$new_n1498)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10430 (
        .A($abc$9276$new_n1489), .B($abc$9276$new_n1498), .Y($abc$9276$new_n1499)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10431 (
        .A($abc$9276$new_n1499), .Y($abc$9276$new_n1500)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10432 (
        .A($abc$9276$new_n1437), .B($abc$9276$new_n1500), .Y(out_0)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10433 (
        .A($abc$9276$new_n381), .B($abc$9276$new_n1003), .Y($abc$9276$new_n1502)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10434 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n1439), .X($abc$9276$new_n1503)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10435 (
        .A($abc$9276$new_n421), .B($abc$9276$new_n1503), .Y($abc$9276$new_n1504)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10436 (
        .A($abc$9276$new_n1504), .Y($abc$9276$new_n1505)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10437 (
        .A($abc$9276$new_n417), .B($abc$9276$new_n1504), .X($abc$9276$new_n1506)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10438 (
        .A(in_35), .B($abc$9276$new_n1502), .Y($abc$9276$new_n1507)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10439 (
        .A($abc$9276$new_n1506), .B($abc$9276$new_n1507), .X($abc$9276$new_n1508)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10440 (
        .A($abc$9276$new_n1508), .Y($abc$9276$new_n1509)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10441 (
        .A(out_0), .B($abc$9276$new_n1509), .Y($abc$9276$new_n1510)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10442 (
        .A(CPU.ABL), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1511)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10443 (
        .A($abc$9276$new_n1510), .B($abc$9276$new_n1511), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8995)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10444 (
        .A($abc$9276$new_n346), .B($abc$9276$new_n449), .Y($abc$9276$new_n1513)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10445 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n449), .X($abc$9276$new_n1514)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10446 (
        .A($abc$9276$new_n1513), .B($abc$9276$new_n1514), .Y($abc$9276$new_n1515)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10447 (
        .A($abc$9276$new_n466), .B($abc$9276$new_n1515), .Y($abc$9276$new_n1516)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10448 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n658), .X($abc$9276$new_n1517)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10449 (
        .A($abc$9276$new_n1517), .Y($abc$9276$new_n1518)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10450 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n684), .X($abc$9276$new_n1519)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10451 (
        .A($abc$9276$new_n1516), .B($abc$9276$new_n1519), .Y($abc$9276$new_n1520)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10452 (
        .A($abc$9276$new_n1518), .B($abc$9276$new_n1520), .X($abc$9276$new_n1521)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10453 (
        .A($abc$9276$new_n407), .B($abc$9276$new_n1521), .X($abc$9276$new_n1522)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10454 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1523)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10455 (
        .A(CPU.ADD), .B($abc$9276$new_n1469), .Y($abc$9276$new_n1524)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10456 (
        .A(CPU.ABL), .B($abc$9276$new_n1480), .Y($abc$9276$new_n1525)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10457 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1483), .Y($abc$9276$new_n1526)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10458 (
        .A($abc$9276$new_n1525), .B($abc$9276$new_n1526), .Y($abc$9276$new_n1527)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10459 (
        .A($abc$9276$new_n1523), .B($abc$9276$new_n1524), .Y($abc$9276$new_n1528)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10460 (
        .A($abc$9276$new_n1043), .B($abc$9276$new_n1528), .X($abc$9276$new_n1529)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10461 (
        .A($abc$9276$new_n1527), .B($abc$9276$new_n1529), .X($abc$9276$new_n1530)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10462 (
        .A($abc$9276$new_n1530), .Y($abc$9276$new_n1531)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10463 (
        .A($abc$9276$new_n1522), .B($abc$9276$new_n1531), .Y(out_1)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10464 (
        .A($abc$9276$new_n1509), .B(out_1), .Y($abc$9276$new_n1533)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10465 (
        .A(CPU.ABL), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1534)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10466 (
        .A($abc$9276$new_n1533), .B($abc$9276$new_n1534), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8997)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10467 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n450), .Y($abc$9276$new_n1536)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10468 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n449), .Y($abc$9276$new_n1537)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10469 (
        .A($abc$9276$new_n1536), .B($abc$9276$new_n1537), .Y($abc$9276$new_n1538)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10470 (
        .A($abc$9276$new_n467), .B($abc$9276$new_n1538), .X($abc$9276$new_n1539)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10471 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n658), .X($abc$9276$new_n1540)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10472 (
        .A($abc$9276$new_n1540), .Y($abc$9276$new_n1541)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10473 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n684), .X($abc$9276$new_n1542)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10474 (
        .A($abc$9276$new_n1539), .B($abc$9276$new_n1542), .Y($abc$9276$new_n1543)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10475 (
        .A($abc$9276$new_n1541), .B($abc$9276$new_n1543), .X($abc$9276$new_n1544)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10476 (
        .A($abc$9276$new_n407), .B($abc$9276$new_n1544), .X($abc$9276$new_n1545)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10477 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1546)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10478 (
        .A(CPU.ADD), .B($abc$9276$new_n1469), .Y($abc$9276$new_n1547)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10479 (
        .A(CPU.ABL), .B($abc$9276$new_n1480), .Y($abc$9276$new_n1548)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10480 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1483), .Y($abc$9276$new_n1549)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10481 (
        .A($abc$9276$new_n1548), .B($abc$9276$new_n1549), .Y($abc$9276$new_n1550)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10482 (
        .A($abc$9276$new_n1063), .B($abc$9276$new_n1550), .X($abc$9276$new_n1551)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10483 (
        .A($abc$9276$new_n1551), .Y($abc$9276$new_n1552)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10484 (
        .A($abc$9276$new_n1547), .B($abc$9276$new_n1552), .Y($abc$9276$new_n1553)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10485 (
        .A($abc$9276$new_n1553), .Y($abc$9276$new_n1554)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10486 (
        .A($abc$9276$new_n1546), .B($abc$9276$new_n1554), .Y($abc$9276$new_n1555)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10487 (
        .A($abc$9276$new_n1555), .Y($abc$9276$new_n1556)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10488 (
        .A($abc$9276$new_n1545), .B($abc$9276$new_n1556), .Y(out_2)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10489 (
        .A($abc$9276$new_n1509), .B(out_2), .Y($abc$9276$new_n1558)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10490 (
        .A(CPU.ABL), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1559)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10491 (
        .A($abc$9276$new_n1558), .B($abc$9276$new_n1559), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8999)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10492 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n450), .Y($abc$9276$new_n1561)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10493 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n449), .Y($abc$9276$new_n1562)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10494 (
        .A($abc$9276$new_n1561), .B($abc$9276$new_n1562), .Y($abc$9276$new_n1563)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10495 (
        .A($abc$9276$new_n467), .B($abc$9276$new_n1563), .X($abc$9276$new_n1564)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10496 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n684), .X($abc$9276$new_n1565)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10497 (
        .A($abc$9276$new_n1565), .Y($abc$9276$new_n1566)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10498 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n658), .X($abc$9276$new_n1567)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10499 (
        .A($abc$9276$new_n1564), .B($abc$9276$new_n1567), .Y($abc$9276$new_n1568)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10500 (
        .A($abc$9276$new_n1566), .B($abc$9276$new_n1568), .X($abc$9276$new_n1569)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10501 (
        .A($abc$9276$new_n407), .B($abc$9276$new_n1569), .X($abc$9276$new_n1570)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10502 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1571)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10503 (
        .A(CPU.ADD), .B($abc$9276$new_n1469), .Y($abc$9276$new_n1572)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10504 (
        .A(CPU.ABL), .B($abc$9276$new_n1480), .Y($abc$9276$new_n1573)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10505 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1483), .Y($abc$9276$new_n1574)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10506 (
        .A($abc$9276$new_n1083), .B($abc$9276$new_n1574), .Y($abc$9276$new_n1575)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10507 (
        .A($abc$9276$new_n1575), .Y($abc$9276$new_n1576)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10508 (
        .A($abc$9276$new_n1573), .B($abc$9276$new_n1576), .Y($abc$9276$new_n1577)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10509 (
        .A($abc$9276$new_n1577), .Y($abc$9276$new_n1578)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10510 (
        .A($abc$9276$new_n1572), .B($abc$9276$new_n1578), .Y($abc$9276$new_n1579)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10511 (
        .A($abc$9276$new_n1579), .Y($abc$9276$new_n1580)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10512 (
        .A($abc$9276$new_n1571), .B($abc$9276$new_n1580), .Y($abc$9276$new_n1581)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10513 (
        .A($abc$9276$new_n1581), .Y($abc$9276$new_n1582)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10514 (
        .A($abc$9276$new_n1570), .B($abc$9276$new_n1582), .Y(out_3)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10515 (
        .A(CPU.ABL), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1584)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10516 (
        .A($abc$9276$new_n1509), .B(out_3), .Y($abc$9276$new_n1585)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10517 (
        .A($abc$9276$new_n1584), .B($abc$9276$new_n1585), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9001)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10518 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n450), .Y($abc$9276$new_n1587)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10519 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n449), .Y($abc$9276$new_n1588)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10520 (
        .A($abc$9276$new_n1587), .B($abc$9276$new_n1588), .Y($abc$9276$new_n1589)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10521 (
        .A($abc$9276$new_n467), .B($abc$9276$new_n1589), .X($abc$9276$new_n1590)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10522 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n658), .X($abc$9276$new_n1591)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10523 (
        .A($abc$9276$new_n1591), .Y($abc$9276$new_n1592)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10524 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n684), .X($abc$9276$new_n1593)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10525 (
        .A($abc$9276$new_n1590), .B($abc$9276$new_n1593), .Y($abc$9276$new_n1594)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10526 (
        .A($abc$9276$new_n1592), .B($abc$9276$new_n1594), .X($abc$9276$new_n1595)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10527 (
        .A($abc$9276$new_n407), .B($abc$9276$new_n1595), .X($abc$9276$new_n1596)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10528 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1597)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10529 (
        .A(CPU.ADD), .B($abc$9276$new_n1469), .Y($abc$9276$new_n1598)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10530 (
        .A(CPU.ABL), .B($abc$9276$new_n1480), .Y($abc$9276$new_n1599)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10531 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1483), .Y($abc$9276$new_n1600)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10532 (
        .A($abc$9276$new_n1100), .B($abc$9276$new_n1600), .Y($abc$9276$new_n1601)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10533 (
        .A($abc$9276$new_n1601), .Y($abc$9276$new_n1602)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10534 (
        .A($abc$9276$new_n1599), .B($abc$9276$new_n1602), .Y($abc$9276$new_n1603)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10535 (
        .A($abc$9276$new_n1603), .Y($abc$9276$new_n1604)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10536 (
        .A($abc$9276$new_n1598), .B($abc$9276$new_n1604), .Y($abc$9276$new_n1605)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10537 (
        .A($abc$9276$new_n1605), .Y($abc$9276$new_n1606)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10538 (
        .A($abc$9276$new_n1597), .B($abc$9276$new_n1606), .Y($abc$9276$new_n1607)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10539 (
        .A($abc$9276$new_n1607), .Y($abc$9276$new_n1608)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10540 (
        .A($abc$9276$new_n1596), .B($abc$9276$new_n1608), .Y(out_4)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10541 (
        .A($abc$9276$new_n1509), .B(out_4), .Y($abc$9276$new_n1610)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10542 (
        .A(CPU.ABL), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1611)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10543 (
        .A($abc$9276$new_n1610), .B($abc$9276$new_n1611), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9003)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10544 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n450), .Y($abc$9276$new_n1613)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10545 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n449), .Y($abc$9276$new_n1614)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10546 (
        .A($abc$9276$new_n1613), .B($abc$9276$new_n1614), .Y($abc$9276$new_n1615)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10547 (
        .A($abc$9276$new_n467), .B($abc$9276$new_n1615), .X($abc$9276$new_n1616)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10548 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n658), .X($abc$9276$new_n1617)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10549 (
        .A($abc$9276$new_n1617), .Y($abc$9276$new_n1618)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10550 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n684), .X($abc$9276$new_n1619)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10551 (
        .A($abc$9276$new_n1616), .B($abc$9276$new_n1619), .Y($abc$9276$new_n1620)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10552 (
        .A($abc$9276$new_n1618), .B($abc$9276$new_n1620), .X($abc$9276$new_n1621)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10553 (
        .A($abc$9276$new_n407), .B($abc$9276$new_n1621), .X($abc$9276$new_n1622)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10554 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1623)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10555 (
        .A(CPU.ADD), .B($abc$9276$new_n1469), .Y($abc$9276$new_n1624)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10556 (
        .A(CPU.ABL), .B($abc$9276$new_n1480), .Y($abc$9276$new_n1625)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10557 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1483), .Y($abc$9276$new_n1626)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10558 (
        .A($abc$9276$new_n1117), .B($abc$9276$new_n1626), .Y($abc$9276$new_n1627)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10559 (
        .A($abc$9276$new_n1627), .Y($abc$9276$new_n1628)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10560 (
        .A($abc$9276$new_n1625), .B($abc$9276$new_n1628), .Y($abc$9276$new_n1629)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10561 (
        .A($abc$9276$new_n1629), .Y($abc$9276$new_n1630)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10562 (
        .A($abc$9276$new_n1624), .B($abc$9276$new_n1630), .Y($abc$9276$new_n1631)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10563 (
        .A($abc$9276$new_n1631), .Y($abc$9276$new_n1632)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10564 (
        .A($abc$9276$new_n1623), .B($abc$9276$new_n1632), .Y($abc$9276$new_n1633)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10565 (
        .A($abc$9276$new_n1633), .Y($abc$9276$new_n1634)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10566 (
        .A($abc$9276$new_n1622), .B($abc$9276$new_n1634), .Y(out_5)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10567 (
        .A($abc$9276$new_n1509), .B(out_5), .Y($abc$9276$new_n1636)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10568 (
        .A(CPU.ABL), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1637)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10569 (
        .A($abc$9276$new_n1636), .B($abc$9276$new_n1637), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9005)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10570 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n450), .Y($abc$9276$new_n1639)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10571 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n449), .Y($abc$9276$new_n1640)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10572 (
        .A($abc$9276$new_n1639), .B($abc$9276$new_n1640), .Y($abc$9276$new_n1641)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10573 (
        .A($abc$9276$new_n467), .B($abc$9276$new_n1641), .X($abc$9276$new_n1642)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10574 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n658), .X($abc$9276$new_n1643)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10575 (
        .A($abc$9276$new_n1643), .Y($abc$9276$new_n1644)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10576 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n684), .X($abc$9276$new_n1645)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10577 (
        .A($abc$9276$new_n1642), .B($abc$9276$new_n1645), .Y($abc$9276$new_n1646)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10578 (
        .A($abc$9276$new_n1644), .B($abc$9276$new_n1646), .X($abc$9276$new_n1647)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10579 (
        .A($abc$9276$new_n407), .B($abc$9276$new_n1647), .X($abc$9276$new_n1648)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10580 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1649)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10581 (
        .A(CPU.ADD), .B($abc$9276$new_n1469), .Y($abc$9276$new_n1650)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10582 (
        .A(CPU.ABL), .B($abc$9276$new_n1480), .Y($abc$9276$new_n1651)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10583 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1483), .Y($abc$9276$new_n1652)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10584 (
        .A($abc$9276$new_n1135), .B($abc$9276$new_n1652), .Y($abc$9276$new_n1653)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10585 (
        .A($abc$9276$new_n1653), .Y($abc$9276$new_n1654)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10586 (
        .A($abc$9276$new_n1651), .B($abc$9276$new_n1654), .Y($abc$9276$new_n1655)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10587 (
        .A($abc$9276$new_n1655), .Y($abc$9276$new_n1656)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10588 (
        .A($abc$9276$new_n1650), .B($abc$9276$new_n1656), .Y($abc$9276$new_n1657)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10589 (
        .A($abc$9276$new_n1657), .Y($abc$9276$new_n1658)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10590 (
        .A($abc$9276$new_n1649), .B($abc$9276$new_n1658), .Y($abc$9276$new_n1659)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10591 (
        .A($abc$9276$new_n1659), .Y($abc$9276$new_n1660)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10592 (
        .A($abc$9276$new_n1648), .B($abc$9276$new_n1660), .Y(out_6)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10593 (
        .A(CPU.ABL), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1662)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10594 (
        .A($abc$9276$new_n1509), .B(out_6), .Y($abc$9276$new_n1663)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10595 (
        .A($abc$9276$new_n1662), .B($abc$9276$new_n1663), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9007)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10596 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n450), .Y($abc$9276$new_n1665)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10597 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n449), .Y($abc$9276$new_n1666)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10598 (
        .A($abc$9276$new_n1665), .B($abc$9276$new_n1666), .Y($abc$9276$new_n1667)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10599 (
        .A($abc$9276$new_n467), .B($abc$9276$new_n1667), .X($abc$9276$new_n1668)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10600 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n684), .X($abc$9276$new_n1669)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10601 (
        .A($abc$9276$new_n1669), .Y($abc$9276$new_n1670)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10602 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n658), .X($abc$9276$new_n1671)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10603 (
        .A($abc$9276$new_n1668), .B($abc$9276$new_n1671), .Y($abc$9276$new_n1672)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10604 (
        .A($abc$9276$new_n1670), .B($abc$9276$new_n1672), .X($abc$9276$new_n1673)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10605 (
        .A($abc$9276$new_n407), .B($abc$9276$new_n1673), .X($abc$9276$new_n1674)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10606 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1675)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10607 (
        .A(CPU.ALU.N), .B($abc$9276$new_n1469), .Y($abc$9276$new_n1676)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10608 (
        .A(CPU.ABL), .B($abc$9276$new_n1480), .Y($abc$9276$new_n1677)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10609 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1483), .Y($abc$9276$new_n1678)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10610 (
        .A($abc$9276$new_n1678), .Y($abc$9276$new_n1679)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10611 (
        .A($abc$9276$new_n1152), .B($abc$9276$new_n1674), .Y($abc$9276$new_n1680)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10612 (
        .A($abc$9276$new_n1676), .B($abc$9276$new_n1677), .Y($abc$9276$new_n1681)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10613 (
        .A($abc$9276$new_n1681), .Y($abc$9276$new_n1682)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10614 (
        .A($abc$9276$new_n1675), .B($abc$9276$new_n1682), .Y($abc$9276$new_n1683)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10615 (
        .A($abc$9276$new_n1679), .B($abc$9276$new_n1683), .X($abc$9276$new_n1684)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10616 (
        .A($abc$9276$new_n1680), .B($abc$9276$new_n1684), .X(out_7)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10617 (
        .A($abc$9276$new_n1509), .B(out_7), .Y($abc$9276$new_n1686)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10618 (
        .A(CPU.ABL), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1687)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10619 (
        .A($abc$9276$new_n1686), .B($abc$9276$new_n1687), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9009)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10620 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1689)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10621 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1467), .Y($abc$9276$new_n1690)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10622 (
        .A($abc$9276$new_n1458), .B($abc$9276$new_n1690), .Y($abc$9276$new_n1691)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10623 (
        .A($abc$9276$new_n407), .B($abc$9276$new_n1170), .Y($abc$9276$new_n1692)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10624 (
        .A(CPU.ABH), .B($abc$9276$new_n1479), .Y($abc$9276$new_n1693)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10625 (
        .A(CPU.ADD), .B($abc$9276$new_n1474), .Y($abc$9276$new_n1694)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10626 (
        .A($abc$9276$new_n1693), .B($abc$9276$new_n1694), .Y($abc$9276$new_n1695)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10627 (
        .A($abc$9276$new_n1692), .B($abc$9276$new_n1695), .X($abc$9276$new_n1696)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10628 (
        .A($abc$9276$new_n1691), .B($abc$9276$new_n1696), .X($abc$9276$new_n1697)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10629 (
        .A($abc$9276$new_n1697), .Y($abc$9276$new_n1698)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10630 (
        .A($abc$9276$new_n1689), .B($abc$9276$new_n1698), .Y(out_8)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10631 (
        .A(CPU.ABH), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1700)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10632 (
        .A($abc$9276$new_n1509), .B(out_8), .Y($abc$9276$new_n1701)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10633 (
        .A($abc$9276$new_n1700), .B($abc$9276$new_n1701), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9011)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10634 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1703)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10635 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1467), .Y($abc$9276$new_n1704)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10636 (
        .A(CPU.ABH), .B($abc$9276$new_n1479), .Y($abc$9276$new_n1705)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10637 (
        .A(CPU.ADD), .B($abc$9276$new_n1474), .Y($abc$9276$new_n1706)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10638 (
        .A($abc$9276$new_n1190), .B($abc$9276$new_n1706), .Y($abc$9276$new_n1707)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10639 (
        .A($abc$9276$new_n1704), .B($abc$9276$new_n1705), .Y($abc$9276$new_n1708)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10640 (
        .A($abc$9276$new_n1707), .B($abc$9276$new_n1708), .X($abc$9276$new_n1709)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10641 (
        .A($abc$9276$new_n1709), .Y($abc$9276$new_n1710)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10642 (
        .A($abc$9276$new_n1703), .B($abc$9276$new_n1710), .Y(out_9)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10643 (
        .A(CPU.ABH), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1712)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10644 (
        .A($abc$9276$new_n1509), .B(out_9), .Y($abc$9276$new_n1713)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10645 (
        .A($abc$9276$new_n1712), .B($abc$9276$new_n1713), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9013)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10646 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1715)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10647 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1467), .Y($abc$9276$new_n1716)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10648 (
        .A(CPU.ADD), .B($abc$9276$new_n1474), .Y($abc$9276$new_n1717)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10649 (
        .A(CPU.ABH), .B($abc$9276$new_n1479), .Y($abc$9276$new_n1718)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10650 (
        .A($abc$9276$new_n1716), .B($abc$9276$new_n1718), .Y($abc$9276$new_n1719)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10651 (
        .A($abc$9276$new_n1210), .B($abc$9276$new_n1717), .Y($abc$9276$new_n1720)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10652 (
        .A($abc$9276$new_n1719), .B($abc$9276$new_n1720), .X($abc$9276$new_n1721)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10653 (
        .A($abc$9276$new_n1721), .Y($abc$9276$new_n1722)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10654 (
        .A($abc$9276$new_n1715), .B($abc$9276$new_n1722), .Y(out_10)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10655 (
        .A(CPU.ABH), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1724)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10656 (
        .A($abc$9276$new_n1509), .B(out_10), .Y($abc$9276$new_n1725)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10657 (
        .A($abc$9276$new_n1724), .B($abc$9276$new_n1725), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9015)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10658 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1727)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10659 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1467), .Y($abc$9276$new_n1728)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10660 (
        .A(CPU.ADD), .B($abc$9276$new_n1474), .Y($abc$9276$new_n1729)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10661 (
        .A(CPU.ABH), .B($abc$9276$new_n1479), .Y($abc$9276$new_n1730)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10662 (
        .A($abc$9276$new_n1230), .B($abc$9276$new_n1730), .Y($abc$9276$new_n1731)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10663 (
        .A($abc$9276$new_n1728), .B($abc$9276$new_n1729), .Y($abc$9276$new_n1732)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10664 (
        .A($abc$9276$new_n1731), .B($abc$9276$new_n1732), .X($abc$9276$new_n1733)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10665 (
        .A($abc$9276$new_n1733), .Y($abc$9276$new_n1734)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10666 (
        .A($abc$9276$new_n1727), .B($abc$9276$new_n1734), .Y(out_11)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10667 (
        .A($abc$9276$new_n1509), .B(out_11), .Y($abc$9276$new_n1736)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10668 (
        .A(CPU.ABH), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1737)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10669 (
        .A($abc$9276$new_n1736), .B($abc$9276$new_n1737), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9017)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10670 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1739)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10671 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1467), .Y($abc$9276$new_n1740)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10672 (
        .A(CPU.ADD), .B($abc$9276$new_n1474), .Y($abc$9276$new_n1741)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10673 (
        .A(CPU.ABH), .B($abc$9276$new_n1479), .Y($abc$9276$new_n1742)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10674 (
        .A($abc$9276$new_n1740), .B($abc$9276$new_n1742), .Y($abc$9276$new_n1743)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10675 (
        .A($abc$9276$new_n1251), .B($abc$9276$new_n1741), .Y($abc$9276$new_n1744)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10676 (
        .A($abc$9276$new_n1743), .B($abc$9276$new_n1744), .X($abc$9276$new_n1745)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10677 (
        .A($abc$9276$new_n1745), .Y($abc$9276$new_n1746)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10678 (
        .A($abc$9276$new_n1739), .B($abc$9276$new_n1746), .Y(out_12)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10679 (
        .A($abc$9276$new_n1509), .B(out_12), .Y($abc$9276$new_n1748)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10680 (
        .A(CPU.ABH), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1749)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10681 (
        .A($abc$9276$new_n1748), .B($abc$9276$new_n1749), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9019)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10682 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1751)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10683 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1467), .Y($abc$9276$new_n1752)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10684 (
        .A(CPU.ABH), .B($abc$9276$new_n1479), .Y($abc$9276$new_n1753)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10685 (
        .A(CPU.ADD), .B($abc$9276$new_n1474), .Y($abc$9276$new_n1754)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10686 (
        .A($abc$9276$new_n1270), .B($abc$9276$new_n1754), .Y($abc$9276$new_n1755)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10687 (
        .A($abc$9276$new_n1752), .B($abc$9276$new_n1753), .Y($abc$9276$new_n1756)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10688 (
        .A($abc$9276$new_n1755), .B($abc$9276$new_n1756), .X($abc$9276$new_n1757)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10689 (
        .A($abc$9276$new_n1757), .Y($abc$9276$new_n1758)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10690 (
        .A($abc$9276$new_n1751), .B($abc$9276$new_n1758), .Y(out_13)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10691 (
        .A($abc$9276$new_n1509), .B(out_13), .Y($abc$9276$new_n1760)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10692 (
        .A(CPU.ABH), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1761)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10693 (
        .A($abc$9276$new_n1760), .B($abc$9276$new_n1761), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9021)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10694 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1763)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10695 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1467), .Y($abc$9276$new_n1764)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10696 (
        .A($abc$9276$new_n1764), .Y($abc$9276$new_n1765)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10697 (
        .A(CPU.ADD), .B($abc$9276$new_n1474), .Y($abc$9276$new_n1766)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10698 (
        .A($abc$9276$new_n1766), .Y($abc$9276$new_n1767)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10699 (
        .A(CPU.ABH), .B($abc$9276$new_n1479), .Y($abc$9276$new_n1768)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10700 (
        .A($abc$9276$new_n1288), .B($abc$9276$new_n1768), .Y($abc$9276$new_n1769)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10701 (
        .A($abc$9276$new_n1767), .B($abc$9276$new_n1769), .X($abc$9276$new_n1770)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10702 (
        .A($abc$9276$new_n1765), .B($abc$9276$new_n1770), .X($abc$9276$new_n1771)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10703 (
        .A($abc$9276$new_n1771), .Y($abc$9276$new_n1772)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10704 (
        .A($abc$9276$new_n1763), .B($abc$9276$new_n1772), .Y(out_14)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10705 (
        .A($abc$9276$new_n1509), .B(out_14), .Y($abc$9276$new_n1774)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10706 (
        .A(CPU.ABH), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1775)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10707 (
        .A($abc$9276$new_n1774), .B($abc$9276$new_n1775), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9023)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10708 (
        .A(CPU.PC), .B($abc$9276$new_n1488), .Y($abc$9276$new_n1777)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10709 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1467), .Y($abc$9276$new_n1778)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10710 (
        .A(CPU.ALU.N), .B($abc$9276$new_n1474), .Y($abc$9276$new_n1779)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10711 (
        .A(CPU.ABH), .B($abc$9276$new_n1479), .Y($abc$9276$new_n1780)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10712 (
        .A($abc$9276$new_n1308), .B($abc$9276$new_n1780), .Y($abc$9276$new_n1781)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10713 (
        .A($abc$9276$new_n1778), .B($abc$9276$new_n1779), .Y($abc$9276$new_n1782)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10714 (
        .A($abc$9276$new_n1781), .B($abc$9276$new_n1782), .X($abc$9276$new_n1783)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10715 (
        .A($abc$9276$new_n1783), .Y($abc$9276$new_n1784)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10716 (
        .A($abc$9276$new_n1777), .B($abc$9276$new_n1784), .Y(out_15)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10717 (
        .A($abc$9276$new_n1509), .B(out_15), .Y($abc$9276$new_n1786)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10718 (
        .A(CPU.ABH), .B($abc$9276$new_n1508), .Y($abc$9276$new_n1787)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10719 (
        .A($abc$9276$new_n1786), .B($abc$9276$new_n1787), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9025)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10720 (
        .A(in_35), .B($abc$9276$new_n1504), .Y($abc$9276$new_n1789)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10721 (
        .A($abc$9276$new_n378), .B($abc$9276$new_n1789), .X($abc$9276$new_n1790)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10722 (
        .A($abc$9276$new_n1790), .Y($abc$9276$new_n1791)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10723 (
        .A($abc$9276$new_n487), .B($abc$9276$new_n1790), .X($abc$9276$new_n1792)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10724 (
        .A(CPU.IRHOLD), .B($abc$9276$new_n1790), .Y($abc$9276$new_n1793)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10725 (
        .A($abc$9276$new_n1792), .B($abc$9276$new_n1793), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9027)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10726 (
        .A($abc$9276$new_n505), .B($abc$9276$new_n1790), .X($abc$9276$new_n1795)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10727 (
        .A(CPU.IRHOLD), .B($abc$9276$new_n1790), .Y($abc$9276$new_n1796)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10728 (
        .A($abc$9276$new_n1795), .B($abc$9276$new_n1796), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9029)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10729 (
        .A(CPU.IRHOLD), .B($abc$9276$new_n1790), .Y($abc$9276$new_n1798)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10730 (
        .A($abc$9276$new_n525), .B($abc$9276$new_n1790), .X($abc$9276$new_n1799)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10731 (
        .A($abc$9276$new_n1798), .B($abc$9276$new_n1799), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9031)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10732 (
        .A($abc$9276$new_n545), .B($abc$9276$new_n1790), .X($abc$9276$new_n1801)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10733 (
        .A(CPU.IRHOLD), .B($abc$9276$new_n1790), .Y($abc$9276$new_n1802)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10734 (
        .A($abc$9276$new_n1801), .B($abc$9276$new_n1802), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9033)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10735 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1791), .Y($abc$9276$new_n1804)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10736 (
        .A(CPU.IRHOLD), .B($abc$9276$new_n1790), .Y($abc$9276$new_n1805)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10737 (
        .A($abc$9276$new_n1804), .B($abc$9276$new_n1805), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9035)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10738 (
        .A(CPU.IRHOLD), .B($abc$9276$new_n1790), .Y($abc$9276$new_n1807)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10739 (
        .A($abc$9276$new_n586), .B($abc$9276$new_n1790), .X($abc$9276$new_n1808)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10740 (
        .A($abc$9276$new_n1807), .B($abc$9276$new_n1808), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9037)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10741 (
        .A(CPU.IRHOLD), .B($abc$9276$new_n1790), .Y($abc$9276$new_n1810)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10742 (
        .A($abc$9276$new_n606), .B($abc$9276$new_n1790), .X($abc$9276$new_n1811)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10743 (
        .A($abc$9276$new_n1810), .B($abc$9276$new_n1811), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9039)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10744 (
        .A(CPU.IRHOLD), .B($abc$9276$new_n1790), .Y($abc$9276$new_n1813)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10745 (
        .A(CPU.DIMUX), .B($abc$9276$new_n1791), .Y($abc$9276$new_n1814)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10746 (
        .A($abc$9276$new_n1813), .B($abc$9276$new_n1814), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9041)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10747 (
        .A($abc$9276$new_n790), .B($abc$9276$new_n882), .Y($abc$9276$new_n1816)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10748 (
        .A($abc$9276$new_n881), .B($abc$9276$new_n1816), .Y($abc$9276$new_n1817)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10749 (
        .A($abc$9276$new_n1817), .Y($abc$9276$new_n1818)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10750 (
        .A($abc$9276$new_n788), .B($abc$9276$new_n816), .X($abc$9276$new_n1819)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10751 (
        .A($abc$9276$new_n787), .B($abc$9276$new_n846), .X($abc$9276$new_n1820)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10752 (
        .A($abc$9276$new_n880), .B($abc$9276$new_n1820), .X($abc$9276$new_n1821)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10753 (
        .A($abc$9276$new_n1819), .B($abc$9276$new_n1821), .Y($abc$9276$new_n1822)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10754 (
        .A($abc$9276$new_n803), .B($abc$9276$new_n932), .X($abc$9276$new_n1823)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10755 (
        .A($abc$9276$new_n778), .B($abc$9276$new_n1823), .X($abc$9276$new_n1824)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10756 (
        .A($abc$9276$new_n1824), .Y($abc$9276$new_n1825)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10757 (
        .A($abc$9276$new_n813), .B($abc$9276$new_n878), .X($abc$9276$new_n1826)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10758 (
        .A($abc$9276$new_n933), .B($abc$9276$new_n1826), .Y($abc$9276$new_n1827)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10759 (
        .A($abc$9276$new_n428), .B($abc$9276$new_n1827), .X($abc$9276$new_n1828)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10760 (
        .A($abc$9276$new_n1825), .B($abc$9276$new_n1828), .X($abc$9276$new_n1829)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10761 (
        .A($abc$9276$new_n814), .B($abc$9276$new_n878), .Y($abc$9276$new_n1830)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10762 (
        .A($abc$9276$new_n1830), .Y($abc$9276$new_n1831)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10763 (
        .A($abc$9276$new_n864), .B($abc$9276$new_n889), .Y($abc$9276$new_n1832)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10764 (
        .A($abc$9276$new_n1831), .B($abc$9276$new_n1832), .Y($abc$9276$new_n1833)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10765 (
        .A($abc$9276$new_n816), .B($abc$9276$new_n821), .X($abc$9276$new_n1834)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10766 (
        .A($abc$9276$new_n1834), .Y($abc$9276$new_n1835)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10767 (
        .A($abc$9276$new_n1833), .B($abc$9276$new_n1834), .Y($abc$9276$new_n1836)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10768 (
        .A($abc$9276$new_n1829), .B($abc$9276$new_n1836), .X($abc$9276$new_n1837)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10769 (
        .A($abc$9276$new_n1822), .B($abc$9276$new_n1837), .X($abc$9276$new_n1838)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10770 (
        .A($abc$9276$new_n1818), .B($abc$9276$new_n1838), .X($abc$9276$new_n1839)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10771 (
        .A($abc$9276$new_n782), .B($abc$9276$new_n816), .X($abc$9276$new_n1840)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10772 (
        .A($abc$9276$new_n865), .B($abc$9276$new_n1840), .Y($abc$9276$new_n1841)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10773 (
        .A($abc$9276$new_n781), .B($abc$9276$new_n890), .X($abc$9276$new_n1842)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10774 (
        .A($abc$9276$new_n1823), .B($abc$9276$new_n1842), .X($abc$9276$new_n1843)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10775 (
        .A($abc$9276$new_n880), .B($abc$9276$new_n1842), .X($abc$9276$new_n1844)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10776 (
        .A($abc$9276$new_n1843), .B($abc$9276$new_n1844), .Y($abc$9276$new_n1845)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10777 (
        .A($abc$9276$new_n1841), .B($abc$9276$new_n1845), .X($abc$9276$new_n1846)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10778 (
        .A($abc$9276$new_n777), .B($abc$9276$new_n935), .X($abc$9276$new_n1847)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10779 (
        .A($abc$9276$new_n801), .B($abc$9276$new_n882), .X($abc$9276$new_n1848)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10780 (
        .A($abc$9276$new_n932), .B($abc$9276$new_n1848), .X($abc$9276$new_n1849)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10781 (
        .A($abc$9276$new_n1847), .B($abc$9276$new_n1849), .Y($abc$9276$new_n1850)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10782 (
        .A($abc$9276$new_n822), .B($abc$9276$new_n1823), .X($abc$9276$new_n1851)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10783 (
        .A($abc$9276$new_n935), .B($abc$9276$new_n1830), .Y($abc$9276$new_n1852)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10784 (
        .A($abc$9276$new_n777), .B($abc$9276$new_n1852), .Y($abc$9276$new_n1853)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10785 (
        .A($abc$9276$new_n788), .B($abc$9276$new_n1823), .X($abc$9276$new_n1854)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10786 (
        .A($abc$9276$new_n1853), .B($abc$9276$new_n1854), .Y($abc$9276$new_n1855)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10787 (
        .A($abc$9276$new_n1855), .Y($abc$9276$new_n1856)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10788 (
        .A($abc$9276$new_n1851), .B($abc$9276$new_n1856), .Y($abc$9276$new_n1857)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10789 (
        .A($abc$9276$new_n1850), .B($abc$9276$new_n1857), .X($abc$9276$new_n1858)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10790 (
        .A($abc$9276$new_n1846), .B($abc$9276$new_n1858), .X($abc$9276$new_n1859)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10791 (
        .A($abc$9276$new_n1839), .B($abc$9276$new_n1859), .X($abc$9276$new_n1860)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10792 (
        .A($abc$9276$new_n985), .B($abc$9276$new_n1502), .Y($abc$9276$new_n1861)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10793 (
        .A($abc$9276$new_n736), .B($abc$9276$new_n1475), .Y($abc$9276$new_n1862)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10794 (
        .A($abc$9276$new_n997), .B($abc$9276$new_n1862), .X($abc$9276$new_n1863)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10795 (
        .A($abc$9276$new_n1861), .B($abc$9276$new_n1863), .X($abc$9276$new_n1864)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10796 (
        .A($abc$9276$new_n1463), .B($abc$9276$new_n1470), .Y($abc$9276$new_n1865)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10797 (
        .A($abc$9276$new_n1010), .B($abc$9276$new_n1865), .X($abc$9276$new_n1866)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10798 (
        .A($abc$9276$new_n1352), .B($abc$9276$new_n1866), .X($abc$9276$new_n1867)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10799 (
        .A($abc$9276$new_n1867), .Y($abc$9276$new_n1868)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10800 (
        .A($abc$9276$new_n389), .B($abc$9276$new_n1003), .Y($abc$9276$new_n1869)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10801 (
        .A($abc$9276$new_n410), .B($abc$9276$new_n998), .Y($abc$9276$new_n1870)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10802 (
        .A($abc$9276$new_n1870), .Y($abc$9276$new_n1871)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10803 (
        .A($abc$9276$new_n1869), .B($abc$9276$new_n1871), .Y($abc$9276$new_n1872)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10804 (
        .A($abc$9276$new_n435), .B($abc$9276$new_n437), .Y($abc$9276$new_n1873)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10805 (
        .A($abc$9276$new_n402), .B($abc$9276$new_n433), .Y($abc$9276$new_n1874)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10806 (
        .A($abc$9276$new_n1873), .B($abc$9276$new_n1874), .X($abc$9276$new_n1875)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10807 (
        .A($abc$9276$new_n1872), .B($abc$9276$new_n1875), .X($abc$9276$new_n1876)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10808 (
        .A($abc$9276$new_n1867), .B($abc$9276$new_n1876), .X($abc$9276$new_n1877)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10809 (
        .A($abc$9276$new_n1864), .B($abc$9276$new_n1877), .X($abc$9276$new_n1878)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10810 (
        .A($abc$9276$new_n729), .B($abc$9276$new_n1446), .Y($abc$9276$new_n1879)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10811 (
        .A($abc$9276$new_n1452), .B($abc$9276$new_n1879), .X($abc$9276$new_n1880)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10812 (
        .A($abc$9276$new_n1015), .B($abc$9276$new_n1880), .X($abc$9276$new_n1881)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10813 (
        .A($abc$9276$new_n453), .B($abc$9276$new_n1005), .X($abc$9276$new_n1882)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10814 (
        .A($abc$9276$new_n1881), .B($abc$9276$new_n1882), .X($abc$9276$new_n1883)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10815 (
        .A($abc$9276$new_n1462), .B($abc$9276$new_n1504), .X($abc$9276$new_n1884)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10816 (
        .A($abc$9276$new_n1464), .B($abc$9276$new_n1472), .Y($abc$9276$new_n1885)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10817 (
        .A($abc$9276$new_n1447), .B($abc$9276$new_n1453), .Y($abc$9276$new_n1886)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10818 (
        .A($abc$9276$new_n1885), .B($abc$9276$new_n1886), .X($abc$9276$new_n1887)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10819 (
        .A($abc$9276$new_n1884), .B($abc$9276$new_n1887), .X($abc$9276$new_n1888)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10820 (
        .A($abc$9276$new_n1477), .B($abc$9276$new_n1482), .Y($abc$9276$new_n1889)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10821 (
        .A($abc$9276$new_n388), .B($abc$9276$new_n396), .X($abc$9276$new_n1890)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10822 (
        .A($abc$9276$new_n1890), .Y($abc$9276$new_n1891)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10823 (
        .A($abc$9276$new_n388), .B($abc$9276$new_n976), .X($abc$9276$new_n1892)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10824 (
        .A($abc$9276$new_n1892), .Y($abc$9276$new_n1893)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10825 (
        .A($abc$9276$new_n1890), .B($abc$9276$new_n1892), .Y($abc$9276$new_n1894)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10826 (
        .A($abc$9276$new_n1889), .B($abc$9276$new_n1894), .X($abc$9276$new_n1895)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10827 (
        .A($abc$9276$new_n397), .B($abc$9276$new_n398), .Y($abc$9276$new_n1896)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10828 (
        .A($abc$9276$new_n1441), .B($abc$9276$new_n1896), .X($abc$9276$new_n1897)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10829 (
        .A($abc$9276$new_n1895), .B($abc$9276$new_n1897), .X($abc$9276$new_n1898)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10830 (
        .A($abc$9276$new_n1888), .B($abc$9276$new_n1898), .X($abc$9276$new_n1899)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10831 (
        .A($abc$9276$new_n1883), .B($abc$9276$new_n1899), .X($abc$9276$new_n1900)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10832 (
        .A($abc$9276$new_n1878), .B($abc$9276$new_n1900), .X($abc$9276$new_n1901)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10833 (
        .A(in_35), .B($abc$9276$new_n1901), .Y($abc$9276$new_n1902)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10834 (
        .A($abc$9276$new_n1902), .Y($abc$9276$new_n1903)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10835 (
        .A($abc$9276$new_n1820), .B($abc$9276$new_n1823), .X($abc$9276$new_n1904)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10836 (
        .A($abc$9276$new_n790), .B($abc$9276$new_n1823), .X($abc$9276$new_n1905)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10837 (
        .A($abc$9276$new_n1860), .B($abc$9276$new_n1903), .Y($abc$9276$new_n1906)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10838 (
        .A($abc$9276$new_n1906), .Y($abc$9276$new_n1907)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10839 (
        .A($abc$9276$new_n775), .B($abc$9276$new_n1826), .X($abc$9276$new_n1908)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10840 (
        .A($abc$9276$new_n1908), .Y($abc$9276$new_n1909)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10841 (
        .A($abc$9276$new_n1850), .B($abc$9276$new_n1909), .X($abc$9276$new_n1910)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10842 (
        .A($abc$9276$new_n1825), .B($abc$9276$new_n1910), .X($abc$9276$new_n1911)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10843 (
        .A($abc$9276$new_n1834), .B($abc$9276$new_n1843), .Y($abc$9276$new_n1912)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10844 (
        .A($abc$9276$new_n1911), .B($abc$9276$new_n1912), .X($abc$9276$new_n1913)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10845 (
        .A($abc$9276$new_n429), .B($abc$9276$new_n1913), .Y($abc$9276$new_n1914)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10846 (
        .A($abc$9276$new_n1440), .B($abc$9276$new_n1482), .Y($abc$9276$new_n1915)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10847 (
        .A($abc$9276$new_n1885), .B($abc$9276$new_n1915), .X($abc$9276$new_n1916)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10848 (
        .A($abc$9276$new_n977), .B($abc$9276$new_n981), .X($abc$9276$new_n1917)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10849 (
        .A($abc$9276$new_n1892), .B($abc$9276$new_n1917), .Y($abc$9276$new_n1918)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10850 (
        .A($abc$9276$new_n397), .B($abc$9276$new_n1012), .Y($abc$9276$new_n1919)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10851 (
        .A($abc$9276$new_n398), .B($abc$9276$new_n418), .Y($abc$9276$new_n1920)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10852 (
        .A($abc$9276$new_n1919), .B($abc$9276$new_n1920), .X($abc$9276$new_n1921)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10853 (
        .A($abc$9276$new_n1918), .B($abc$9276$new_n1921), .X($abc$9276$new_n1922)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10854 (
        .A($abc$9276$new_n1916), .B($abc$9276$new_n1922), .X($abc$9276$new_n1923)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10855 (
        .A(CPU.store), .B(CPU.ALU.CO), .X($abc$9276$new_n1924)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10856 (
        .A($abc$9276$new_n1924), .Y($abc$9276$new_n1925)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10857 (
        .A(CPU.write_back), .B($abc$9276$new_n1924), .X($abc$9276$new_n1926)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10858 (
        .A($abc$9276$new_n1459), .B($abc$9276$new_n1926), .X($abc$9276$new_n1927)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10859 (
        .A($abc$9276$new_n1869), .B($abc$9276$new_n1927), .Y($abc$9276$new_n1928)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10860 (
        .A($abc$9276$new_n452), .B($abc$9276$new_n1004), .Y($abc$9276$new_n1929)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10861 (
        .A($abc$9276$new_n1928), .B($abc$9276$new_n1929), .X($abc$9276$new_n1930)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10862 (
        .A($abc$9276$new_n437), .B($abc$9276$new_n1446), .Y($abc$9276$new_n1931)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10863 (
        .A($abc$9276$new_n1891), .B($abc$9276$new_n1931), .X($abc$9276$new_n1932)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10864 (
        .A($abc$9276$new_n413), .B($abc$9276$new_n421), .Y($abc$9276$new_n1933)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10865 (
        .A($abc$9276$new_n433), .B($abc$9276$new_n1461), .Y($abc$9276$new_n1934)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10866 (
        .A($abc$9276$new_n1933), .B($abc$9276$new_n1934), .X($abc$9276$new_n1935)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10867 (
        .A($abc$9276$new_n1932), .B($abc$9276$new_n1935), .X($abc$9276$new_n1936)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10868 (
        .A($abc$9276$new_n1930), .B($abc$9276$new_n1936), .X($abc$9276$new_n1937)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10869 (
        .A($abc$9276$new_n1867), .B($abc$9276$new_n1937), .X($abc$9276$new_n1938)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10870 (
        .A($abc$9276$new_n1923), .B($abc$9276$new_n1938), .X($abc$9276$new_n1939)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10871 (
        .A($abc$9276$new_n1939), .Y($abc$9276$new_n1940)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10872 (
        .A($abc$9276$new_n1914), .B($abc$9276$new_n1940), .Y($abc$9276$new_n1941)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10873 (
        .A($abc$9276$new_n1907), .B($abc$9276$new_n1941), .Y($abc$9276$new_n1942)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10874 (
        .A(CPU.state), .B($abc$9276$new_n1906), .Y($abc$9276$new_n1943)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10875 (
        .A($abc$9276$new_n1942), .B($abc$9276$new_n1943), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9043)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10876 (
        .A($abc$9276$new_n934), .B($abc$9276$new_n1844), .Y($abc$9276$new_n1945)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10877 (
        .A($abc$9276$new_n777), .B($abc$9276$new_n933), .X($abc$9276$new_n1946)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10878 (
        .A($abc$9276$new_n1819), .B($abc$9276$new_n1946), .Y($abc$9276$new_n1947)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10879 (
        .A($abc$9276$new_n1947), .Y($abc$9276$new_n1948)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10880 (
        .A($abc$9276$new_n1855), .B($abc$9276$new_n1909), .X($abc$9276$new_n1949)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10881 (
        .A($abc$9276$new_n1947), .B($abc$9276$new_n1949), .X($abc$9276$new_n1950)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10882 (
        .A($abc$9276$new_n1945), .B($abc$9276$new_n1950), .X($abc$9276$new_n1951)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10883 (
        .A($abc$9276$new_n429), .B($abc$9276$new_n1951), .Y($abc$9276$new_n1952)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10884 (
        .A(CPU.cond_code), .B(CPU.cond_code), .X($abc$9276$new_n1953)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10885 (
        .A($abc$9276$new_n1953), .Y($abc$9276$new_n1954)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10886 (
        .A($flatten\CPU.$procmux$291.B), .B($abc$9276$new_n1954), .Y($abc$9276$new_n1955)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10887 (
        .A(CPU.cond_code), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9182), .X($abc$9276$new_n1956)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10888 (
        .A($abc$9276$new_n1956), .Y($abc$9276$new_n1957)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10889 (
        .A($flatten\CPU.$procmux$291.B), .B($abc$9276$new_n1957), .Y($abc$9276$new_n1958)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10890 (
        .A($abc$9276$new_n1955), .B($abc$9276$new_n1958), .Y($abc$9276$new_n1959)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10891 (
        .A($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9184), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9182), .X($abc$9276$new_n1960)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10892 (
        .A($abc$9276$new_n362), .B($abc$9276$new_n1960), .X($abc$9276$new_n1961)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10893 (
        .A(CPU.cond_code), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9184), .X($abc$9276$new_n1962)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10894 (
        .A($abc$9276$new_n363), .B($abc$9276$new_n1962), .X($abc$9276$new_n1963)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10895 (
        .A($abc$9276$new_n1961), .B($abc$9276$new_n1963), .Y($abc$9276$new_n1964)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10896 (
        .A($abc$9276$new_n1959), .B($abc$9276$new_n1964), .X($abc$9276$new_n1965)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10897 (
        .A($abc$9276$new_n379), .B($abc$9276$new_n1965), .Y($abc$9276$new_n1966)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10898 (
        .A($flatten\CPU.$procmux$291.B), .B($abc$9276$new_n1954), .Y($abc$9276$new_n1967)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10899 (
        .A($flatten\CPU.$procmux$291.B), .B($abc$9276$new_n1957), .Y($abc$9276$new_n1968)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10900 (
        .A($abc$9276$new_n1967), .B($abc$9276$new_n1968), .Y($abc$9276$new_n1969)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10901 (
        .A($abc$9276$new_n349), .B($abc$9276$new_n1960), .X($abc$9276$new_n1970)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10902 (
        .A($abc$9276$new_n361), .B($abc$9276$new_n1962), .X($abc$9276$new_n1971)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10903 (
        .A($abc$9276$new_n1970), .B($abc$9276$new_n1971), .Y($abc$9276$new_n1972)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10904 (
        .A($abc$9276$new_n1969), .B($abc$9276$new_n1972), .X($abc$9276$new_n1973)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10905 (
        .A($abc$9276$new_n360), .B($abc$9276$new_n1973), .Y($abc$9276$new_n1974)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10906 (
        .A($abc$9276$new_n1966), .B($abc$9276$new_n1974), .Y($abc$9276$new_n1975)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10907 (
        .A($abc$9276$new_n1002), .B($abc$9276$new_n1975), .Y($abc$9276$new_n1976)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10908 (
        .A($abc$9276$new_n403), .B($abc$9276$new_n422), .X($abc$9276$new_n1977)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10909 (
        .A($abc$9276$new_n1977), .Y($abc$9276$new_n1978)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10910 (
        .A($abc$9276$new_n1446), .B($abc$9276$new_n1481), .Y($abc$9276$new_n1979)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10911 (
        .A($abc$9276$new_n1454), .B($abc$9276$new_n1979), .X($abc$9276$new_n1980)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10912 (
        .A($abc$9276$new_n1918), .B($abc$9276$new_n1980), .X($abc$9276$new_n1981)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10913 (
        .A($abc$9276$new_n1977), .B($abc$9276$new_n1981), .X($abc$9276$new_n1982)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10914 (
        .A(CPU.write_back), .B($abc$9276$new_n1916), .Y($abc$9276$new_n1983)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10915 (
        .A($abc$9276$new_n1983), .Y($abc$9276$new_n1984)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10916 (
        .A($abc$9276$new_n390), .B($abc$9276$new_n1012), .Y($abc$9276$new_n1985)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10917 (
        .A($abc$9276$new_n439), .B($abc$9276$new_n1985), .X($abc$9276$new_n1986)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10918 (
        .A($abc$9276$new_n1477), .B($abc$9276$new_n1503), .Y($abc$9276$new_n1987)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10919 (
        .A($abc$9276$new_n1870), .B($abc$9276$new_n1987), .X($abc$9276$new_n1988)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10920 (
        .A($abc$9276$new_n1986), .B($abc$9276$new_n1988), .X($abc$9276$new_n1989)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10921 (
        .A($abc$9276$new_n1989), .Y($abc$9276$new_n1990)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10922 (
        .A($abc$9276$new_n1976), .B($abc$9276$new_n1990), .Y($abc$9276$new_n1991)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10923 (
        .A($abc$9276$new_n1982), .B($abc$9276$new_n1991), .X($abc$9276$new_n1992)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10924 (
        .A($abc$9276$new_n1984), .B($abc$9276$new_n1992), .X($abc$9276$new_n1993)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10925 (
        .A($abc$9276$new_n1993), .Y($abc$9276$new_n1994)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10926 (
        .A($abc$9276$new_n1952), .B($abc$9276$new_n1994), .Y($abc$9276$new_n1995)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10927 (
        .A($abc$9276$new_n1906), .B($abc$9276$new_n1995), .X($abc$9276$new_n1996)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10928 (
        .A(CPU.state), .B($abc$9276$new_n1907), .X($abc$9276$new_n1997)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10929 (
        .A($abc$9276$new_n1996), .B($abc$9276$new_n1997), .Y($abc$9276$new_n1998)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10930 (
        .A($abc$9276$new_n1998), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9045)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10931 (
        .A($abc$9276$new_n1911), .B($abc$9276$new_n1947), .X($abc$9276$new_n2000)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10932 (
        .A($abc$9276$new_n1846), .B($abc$9276$new_n2000), .X($abc$9276$new_n2001)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10933 (
        .A($abc$9276$new_n429), .B($abc$9276$new_n2001), .Y($abc$9276$new_n2002)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10934 (
        .A($abc$9276$new_n977), .B($abc$9276$new_n1001), .Y($abc$9276$new_n2003)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10935 (
        .A($abc$9276$new_n1448), .B($abc$9276$new_n2003), .X($abc$9276$new_n2004)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10936 (
        .A($abc$9276$new_n1462), .B($abc$9276$new_n1893), .X($abc$9276$new_n2005)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10937 (
        .A($abc$9276$new_n1452), .B($abc$9276$new_n1870), .X($abc$9276$new_n2006)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10938 (
        .A($abc$9276$new_n2005), .B($abc$9276$new_n2006), .X($abc$9276$new_n2007)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10939 (
        .A($abc$9276$new_n2004), .B($abc$9276$new_n2007), .X($abc$9276$new_n2008)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10940 (
        .A($abc$9276$new_n402), .B($abc$9276$new_n423), .Y($abc$9276$new_n2009)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10941 (
        .A($abc$9276$new_n421), .B($abc$9276$new_n1477), .Y($abc$9276$new_n2010)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10942 (
        .A($abc$9276$new_n2010), .Y($abc$9276$new_n2011)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10943 (
        .A($abc$9276$new_n1873), .B($abc$9276$new_n2010), .X($abc$9276$new_n2012)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10944 (
        .A($abc$9276$new_n2009), .B($abc$9276$new_n2012), .X($abc$9276$new_n2013)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10945 (
        .A($abc$9276$new_n1864), .B($abc$9276$new_n2013), .X($abc$9276$new_n2014)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10946 (
        .A($abc$9276$new_n2008), .B($abc$9276$new_n2014), .X($abc$9276$new_n2015)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10947 (
        .A($flatten\CPU.$procmux$415.B), .B($abc$9276$new_n1916), .Y($abc$9276$new_n2016)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10948 (
        .A($abc$9276$new_n1868), .B($abc$9276$new_n2016), .Y($abc$9276$new_n2017)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10949 (
        .A($abc$9276$new_n2017), .Y($abc$9276$new_n2018)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10950 (
        .A($abc$9276$new_n2002), .B($abc$9276$new_n2018), .Y($abc$9276$new_n2019)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10951 (
        .A($abc$9276$new_n2015), .B($abc$9276$new_n2019), .X($abc$9276$new_n2020)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10952 (
        .A($abc$9276$new_n1907), .B($abc$9276$new_n2020), .Y($abc$9276$new_n2021)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10953 (
        .A(CPU.state), .B($abc$9276$new_n1906), .Y($abc$9276$new_n2022)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10954 (
        .A($abc$9276$new_n2021), .B($abc$9276$new_n2022), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9047)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10955 (
        .A($abc$9276$new_n1821), .B($abc$9276$new_n1854), .Y($abc$9276$new_n2024)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10956 (
        .A($abc$9276$new_n1851), .B($abc$9276$new_n1948), .Y($abc$9276$new_n2025)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10957 (
        .A($abc$9276$new_n2024), .B($abc$9276$new_n2025), .X($abc$9276$new_n2026)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10958 (
        .A($abc$9276$new_n1910), .B($abc$9276$new_n2026), .X($abc$9276$new_n2027)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10959 (
        .A($abc$9276$new_n429), .B($abc$9276$new_n2027), .Y($abc$9276$new_n2028)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10960 (
        .A($abc$9276$new_n1461), .B($abc$9276$new_n1924), .X($abc$9276$new_n2029)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10961 (
        .A($abc$9276$new_n2029), .Y($abc$9276$new_n2030)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10962 (
        .A($abc$9276$new_n1927), .B($abc$9276$new_n2011), .Y($abc$9276$new_n2031)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10963 (
        .A($abc$9276$new_n2030), .B($abc$9276$new_n2031), .X($abc$9276$new_n2032)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10964 (
        .A($abc$9276$new_n1864), .B($abc$9276$new_n2032), .X($abc$9276$new_n2033)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10965 (
        .A($abc$9276$new_n437), .B($abc$9276$new_n729), .Y($abc$9276$new_n2034)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10966 (
        .A($abc$9276$new_n2034), .Y($abc$9276$new_n2035)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10967 (
        .A($abc$9276$new_n982), .B($abc$9276$new_n2035), .Y($abc$9276$new_n2036)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10968 (
        .A($abc$9276$new_n1452), .B($abc$9276$new_n1886), .X($abc$9276$new_n2037)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10969 (
        .A($abc$9276$new_n2036), .B($abc$9276$new_n2037), .X($abc$9276$new_n2038)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10970 (
        .A($abc$9276$new_n451), .B($abc$9276$new_n1891), .X($abc$9276$new_n2039)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10971 (
        .A($abc$9276$new_n1921), .B($abc$9276$new_n2039), .X($abc$9276$new_n2040)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10972 (
        .A($abc$9276$new_n2038), .B($abc$9276$new_n2040), .X($abc$9276$new_n2041)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10973 (
        .A($abc$9276$new_n2033), .B($abc$9276$new_n2041), .X($abc$9276$new_n2042)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10974 (
        .A($abc$9276$new_n1001), .B($abc$9276$new_n1975), .X($abc$9276$new_n2043)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10975 (
        .A($abc$9276$new_n2018), .B($abc$9276$new_n2043), .Y($abc$9276$new_n2044)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10976 (
        .A($abc$9276$new_n2042), .B($abc$9276$new_n2044), .X($abc$9276$new_n2045)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10977 (
        .A($abc$9276$new_n2045), .Y($abc$9276$new_n2046)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10978 (
        .A($abc$9276$new_n2028), .B($abc$9276$new_n2046), .Y($abc$9276$new_n2047)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10979 (
        .A($abc$9276$new_n1907), .B($abc$9276$new_n2047), .Y($abc$9276$new_n2048)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10980 (
        .A(CPU.state), .B($abc$9276$new_n1906), .Y($abc$9276$new_n2049)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10981 (
        .A($abc$9276$new_n2048), .B($abc$9276$new_n2049), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9049)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10982 (
        .A($abc$9276$new_n774), .B($abc$9276$new_n1826), .X($abc$9276$new_n2051)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10983 (
        .A($abc$9276$new_n1905), .B($abc$9276$new_n2051), .Y($abc$9276$new_n2052)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10984 (
        .A($abc$9276$new_n1822), .B($abc$9276$new_n2052), .X($abc$9276$new_n2053)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10985 (
        .A($abc$9276$new_n1945), .B($abc$9276$new_n2053), .X($abc$9276$new_n2054)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10986 (
        .A($abc$9276$new_n429), .B($abc$9276$new_n2054), .Y($abc$9276$new_n2055)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10987 (
        .A($abc$9276$new_n1461), .B($abc$9276$new_n1925), .X($abc$9276$new_n2056)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10988 (
        .A($abc$9276$new_n421), .B($abc$9276$new_n1438), .Y($abc$9276$new_n2057)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10989 (
        .A($abc$9276$new_n1447), .B($abc$9276$new_n1892), .Y($abc$9276$new_n2058)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10990 (
        .A($abc$9276$new_n2057), .B($abc$9276$new_n2058), .X($abc$9276$new_n2059)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10991 (
        .A($abc$9276$new_n436), .B($abc$9276$new_n1870), .X($abc$9276$new_n2060)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10992 (
        .A($abc$9276$new_n2059), .B($abc$9276$new_n2060), .X($abc$9276$new_n2061)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10993 (
        .A($abc$9276$new_n2039), .B($abc$9276$new_n2061), .X($abc$9276$new_n2062)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10994 (
        .A($abc$9276$new_n1869), .B($abc$9276$new_n2056), .Y($abc$9276$new_n2063)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10995 (
        .A($abc$9276$new_n2063), .Y($abc$9276$new_n2064)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10996 (
        .A($abc$9276$new_n2055), .B($abc$9276$new_n2064), .Y($abc$9276$new_n2065)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10997 (
        .A($abc$9276$new_n2062), .B($abc$9276$new_n2065), .X($abc$9276$new_n2066)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10998 (
        .A($abc$9276$new_n1907), .B($abc$9276$new_n2066), .Y($abc$9276$new_n2067)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$10999 (
        .A(CPU.state), .B($abc$9276$new_n1906), .Y($abc$9276$new_n2068)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11000 (
        .A($abc$9276$new_n2067), .B($abc$9276$new_n2068), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9051)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11001 (
        .A($abc$9276$new_n1826), .B($abc$9276$new_n1904), .Y($abc$9276$new_n2070)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11002 (
        .A($abc$9276$new_n1841), .B($abc$9276$new_n1912), .X($abc$9276$new_n2071)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11003 (
        .A($abc$9276$new_n2070), .B($abc$9276$new_n2071), .X($abc$9276$new_n2072)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11004 (
        .A($abc$9276$new_n429), .B($abc$9276$new_n2072), .Y($abc$9276$new_n2073)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11005 (
        .A($abc$9276$new_n1874), .B($abc$9276$new_n1920), .X($abc$9276$new_n2074)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11006 (
        .A($abc$9276$new_n417), .B($abc$9276$new_n1987), .X($abc$9276$new_n2075)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11007 (
        .A($abc$9276$new_n1984), .B($abc$9276$new_n2075), .X($abc$9276$new_n2076)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11008 (
        .A($abc$9276$new_n2074), .B($abc$9276$new_n2076), .X($abc$9276$new_n2077)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11009 (
        .A($abc$9276$new_n2077), .Y($abc$9276$new_n2078)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11010 (
        .A($abc$9276$new_n2073), .B($abc$9276$new_n2078), .Y($abc$9276$new_n2079)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11011 (
        .A($abc$9276$new_n1880), .B($abc$9276$new_n2079), .X($abc$9276$new_n2080)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11012 (
        .A($abc$9276$new_n1907), .B($abc$9276$new_n2080), .Y($abc$9276$new_n2081)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11013 (
        .A(CPU.state), .B($abc$9276$new_n1906), .Y($abc$9276$new_n2082)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11014 (
        .A($abc$9276$new_n2081), .B($abc$9276$new_n2082), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9053)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11015 (
        .A(CPU.dst_reg), .B($abc$9276$new_n753), .X($abc$9276$new_n2084)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11016 (
        .A($abc$9276$new_n816), .B($abc$9276$new_n957), .X($abc$9276$new_n2085)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11017 (
        .A($abc$9276$new_n774), .B($abc$9276$new_n814), .X($abc$9276$new_n2086)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11018 (
        .A($abc$9276$new_n2086), .Y($abc$9276$new_n2087)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11019 (
        .A($abc$9276$new_n787), .B($abc$9276$new_n885), .X($abc$9276$new_n2088)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11020 (
        .A($abc$9276$new_n815), .B($abc$9276$new_n2088), .X($abc$9276$new_n2089)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11021 (
        .A($abc$9276$new_n864), .B($abc$9276$new_n918), .X($abc$9276$new_n2090)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11022 (
        .A($abc$9276$new_n803), .B($abc$9276$new_n918), .X($abc$9276$new_n2091)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11023 (
        .A($abc$9276$new_n2087), .B($abc$9276$new_n2091), .X($abc$9276$new_n2092)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11024 (
        .A($abc$9276$new_n2085), .B($abc$9276$new_n2092), .Y($abc$9276$new_n2093)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11025 (
        .A($abc$9276$new_n2089), .B($abc$9276$new_n2090), .Y($abc$9276$new_n2094)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11026 (
        .A($abc$9276$new_n2093), .B($abc$9276$new_n2094), .X($abc$9276$new_n2095)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11027 (
        .A($abc$9276$new_n752), .B($abc$9276$new_n2095), .X($abc$9276$new_n2096)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11028 (
        .A($abc$9276$new_n960), .B($abc$9276$new_n2096), .X($abc$9276$new_n2097)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11029 (
        .A($abc$9276$new_n2084), .B($abc$9276$new_n2097), .Y($abc$9276$new_n2098)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11030 (
        .A($abc$9276$new_n2098), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9057)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11031 (
        .A(CPU.dst_reg), .B($abc$9276$new_n753), .X($abc$9276$new_n2100)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11032 (
        .A($abc$9276$new_n829), .B($abc$9276$new_n853), .X($abc$9276$new_n2101)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11033 (
        .A($abc$9276$new_n865), .B($abc$9276$new_n2101), .X($abc$9276$new_n2102)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11034 (
        .A($abc$9276$new_n2102), .Y($abc$9276$new_n2103)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11035 (
        .A($abc$9276$new_n1835), .B($abc$9276$new_n2093), .X($abc$9276$new_n2104)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11036 (
        .A($abc$9276$new_n2103), .B($abc$9276$new_n2104), .X($abc$9276$new_n2105)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11037 (
        .A($abc$9276$new_n752), .B($abc$9276$new_n2105), .X($abc$9276$new_n2106)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11038 (
        .A($abc$9276$new_n2100), .B($abc$9276$new_n2106), .Y($abc$9276$new_n2107)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11039 (
        .A($abc$9276$new_n2107), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9061)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11040 (
        .A($abc$9276$new_n371), .B($abc$9276$new_n752), .Y($abc$9276$new_n2109)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11041 (
        .A($abc$9276$new_n815), .B($abc$9276$new_n2101), .X($abc$9276$new_n2110)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11042 (
        .A($abc$9276$new_n813), .B($abc$9276$new_n827), .X($abc$9276$new_n2111)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11043 (
        .A($abc$9276$new_n853), .B($abc$9276$new_n2111), .X($abc$9276$new_n2112)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11044 (
        .A($abc$9276$new_n2112), .Y($abc$9276$new_n2113)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11045 (
        .A($abc$9276$new_n958), .B($abc$9276$new_n2110), .Y($abc$9276$new_n2114)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11046 (
        .A($abc$9276$new_n2113), .B($abc$9276$new_n2114), .X($abc$9276$new_n2115)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11047 (
        .A($abc$9276$new_n804), .B($abc$9276$new_n2115), .Y($abc$9276$new_n2116)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11048 (
        .A($abc$9276$new_n753), .B($abc$9276$new_n2085), .Y($abc$9276$new_n2117)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11049 (
        .A($abc$9276$new_n2117), .Y($abc$9276$new_n2118)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11050 (
        .A($abc$9276$new_n2116), .B($abc$9276$new_n2118), .Y($abc$9276$new_n2119)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11051 (
        .A($abc$9276$new_n953), .B($abc$9276$new_n2111), .Y($abc$9276$new_n2120)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11052 (
        .A($abc$9276$new_n938), .B($abc$9276$new_n2120), .Y($abc$9276$new_n2121)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11053 (
        .A($abc$9276$new_n2088), .B($abc$9276$new_n2121), .Y($abc$9276$new_n2122)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11054 (
        .A($abc$9276$new_n960), .B($abc$9276$new_n2122), .X($abc$9276$new_n2123)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11055 (
        .A($abc$9276$new_n2119), .B($abc$9276$new_n2123), .X($abc$9276$new_n2124)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11056 (
        .A($abc$9276$new_n2109), .B($abc$9276$new_n2124), .Y($abc$9276$new_n2125)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11057 (
        .A($abc$9276$new_n2125), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9065)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11058 (
        .A($abc$9276$new_n865), .B($abc$9276$new_n951), .X($abc$9276$new_n2127)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11059 (
        .A($abc$9276$new_n2127), .Y($abc$9276$new_n2128)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11060 (
        .A($abc$9276$new_n2119), .B($abc$9276$new_n2128), .X($abc$9276$new_n2129)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11061 (
        .A(CPU.src_reg), .B($abc$9276$new_n753), .X($abc$9276$new_n2130)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11062 (
        .A($abc$9276$new_n2129), .B($abc$9276$new_n2130), .Y($abc$9276$new_n2131)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11063 (
        .A($abc$9276$new_n2131), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9069)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11064 (
        .A(CPU.op), .B($abc$9276$new_n753), .X($abc$9276$new_n2133)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11065 (
        .A($abc$9276$new_n769), .B($abc$9276$new_n903), .Y($abc$9276$new_n2134)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11066 (
        .A($abc$9276$new_n889), .B($abc$9276$new_n2134), .X($abc$9276$new_n2135)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11067 (
        .A($abc$9276$new_n2135), .Y($abc$9276$new_n2136)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11068 (
        .A($abc$9276$new_n826), .B($abc$9276$new_n864), .X($abc$9276$new_n2137)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11069 (
        .A($abc$9276$new_n2137), .Y($abc$9276$new_n2138)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11070 (
        .A($abc$9276$new_n860), .B($abc$9276$new_n874), .Y($abc$9276$new_n2139)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11071 (
        .A($abc$9276$new_n2138), .B($abc$9276$new_n2139), .X($abc$9276$new_n2140)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11072 (
        .A($abc$9276$new_n752), .B($abc$9276$new_n2140), .X($abc$9276$new_n2141)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11073 (
        .A($abc$9276$new_n2136), .B($abc$9276$new_n2139), .X($abc$9276$new_n2142)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11074 (
        .A($abc$9276$new_n2142), .Y($abc$9276$new_n2143)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11075 (
        .A($abc$9276$new_n2136), .B($abc$9276$new_n2141), .X($abc$9276$new_n2144)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11076 (
        .A($abc$9276$new_n2133), .B($abc$9276$new_n2144), .Y($abc$9276$new_n2145)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11077 (
        .A($abc$9276$new_n2145), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9073)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11078 (
        .A($abc$9276$new_n827), .B($abc$9276$new_n911), .X($abc$9276$new_n2147)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11079 (
        .A($abc$9276$new_n2147), .Y($abc$9276$new_n2148)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11080 (
        .A($abc$9276$new_n789), .B($abc$9276$new_n2085), .X($abc$9276$new_n2149)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11081 (
        .A($abc$9276$new_n839), .B($abc$9276$new_n889), .X($abc$9276$new_n2150)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11082 (
        .A($abc$9276$new_n959), .B($abc$9276$new_n2150), .Y($abc$9276$new_n2151)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11083 (
        .A($abc$9276$new_n2151), .Y($abc$9276$new_n2152)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11084 (
        .A($abc$9276$new_n2149), .B($abc$9276$new_n2152), .Y($abc$9276$new_n2153)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11085 (
        .A($abc$9276$new_n2148), .B($abc$9276$new_n2153), .X($abc$9276$new_n2154)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11086 (
        .A($abc$9276$new_n888), .B($abc$9276$new_n2154), .X($abc$9276$new_n2155)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11087 (
        .A($abc$9276$new_n2142), .B($abc$9276$new_n2155), .X($abc$9276$new_n2156)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11088 (
        .A($abc$9276$new_n753), .B($abc$9276$new_n2156), .Y($abc$9276$new_n2157)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11089 (
        .A(CPU.op), .B($abc$9276$new_n752), .Y($abc$9276$new_n2158)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11090 (
        .A($abc$9276$new_n2157), .B($abc$9276$new_n2158), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9077)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11091 (
        .A(CPU.op), .B($abc$9276$new_n753), .X($abc$9276$new_n2160)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11092 (
        .A($abc$9276$new_n2138), .B($abc$9276$new_n2156), .X($abc$9276$new_n2161)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11093 (
        .A($abc$9276$new_n753), .B($abc$9276$new_n2161), .Y($abc$9276$new_n2162)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11094 (
        .A($abc$9276$new_n864), .B($abc$9276$new_n891), .Y($abc$9276$new_n2163)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11095 (
        .A($abc$9276$new_n780), .B($abc$9276$new_n2163), .Y($abc$9276$new_n2164)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11096 (
        .A($abc$9276$new_n2164), .Y($abc$9276$new_n2165)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11097 (
        .A($abc$9276$new_n2155), .B($abc$9276$new_n2165), .X($abc$9276$new_n2166)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11098 (
        .A($abc$9276$new_n2162), .B($abc$9276$new_n2166), .X($abc$9276$new_n2167)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11099 (
        .A($abc$9276$new_n2160), .B($abc$9276$new_n2167), .Y($abc$9276$new_n2168)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11100 (
        .A($abc$9276$new_n2168), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9081)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11101 (
        .A(CPU.op), .B($abc$9276$new_n753), .X($abc$9276$new_n2170)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11102 (
        .A($abc$9276$new_n786), .B($abc$9276$new_n2135), .X($abc$9276$new_n2171)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11103 (
        .A($abc$9276$new_n2171), .Y($abc$9276$new_n2172)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11104 (
        .A($abc$9276$new_n2141), .B($abc$9276$new_n2172), .X($abc$9276$new_n2173)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11105 (
        .A($abc$9276$new_n2143), .B($abc$9276$new_n2173), .X($abc$9276$new_n2174)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11106 (
        .A($abc$9276$new_n2170), .B($abc$9276$new_n2174), .Y($abc$9276$new_n2175)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11107 (
        .A($abc$9276$new_n2175), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9085)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11108 (
        .A($abc$9276$new_n359), .B(CPU.ALU.BI7), .Y($abc$9276$new_n2177)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11109 (
        .A($abc$9276$new_n978), .B($abc$9276$new_n1462), .X($abc$9276$new_n2178)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11110 (
        .A($abc$9276$new_n428), .B($abc$9276$new_n1464), .Y($abc$9276$new_n2179)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11111 (
        .A($abc$9276$new_n737), .B($abc$9276$new_n1478), .X($abc$9276$new_n2180)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11112 (
        .A($abc$9276$new_n377), .B($abc$9276$new_n2180), .X($abc$9276$new_n2181)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11113 (
        .A($abc$9276$new_n2179), .B($abc$9276$new_n2181), .X($abc$9276$new_n2182)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11114 (
        .A($abc$9276$new_n2178), .B($abc$9276$new_n2182), .X($abc$9276$new_n2183)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11115 (
        .A($abc$9276$new_n2183), .Y($abc$9276$new_n2184)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11116 (
        .A(CPU.rotate), .B(CPU.C), .Y($abc$9276$new_n2185)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11117 (
        .A(CPU.shift), .B(CPU.load_only), .X($abc$9276$new_n2186)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11118 (
        .A(oeb_0), .B($abc$9276$new_n2186), .Y($abc$9276$new_n2187)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11119 (
        .A($abc$9276$new_n363), .B($abc$9276$new_n2186), .X($abc$9276$new_n2188)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11120 (
        .A($abc$9276$new_n2187), .B($abc$9276$new_n2188), .Y($abc$9276$new_n2189)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11121 (
        .A(CPU.compare), .B($abc$9276$new_n2189), .X($abc$9276$new_n2190)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11122 (
        .A($abc$9276$new_n351), .B(CPU.compare), .Y($abc$9276$new_n2191)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11123 (
        .A($abc$9276$new_n2190), .B($abc$9276$new_n2191), .Y($abc$9276$new_n2192)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11124 (
        .A(CPU.rotate), .B($abc$9276$new_n2192), .X($abc$9276$new_n2193)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11125 (
        .A($abc$9276$new_n2185), .B($abc$9276$new_n2193), .Y($abc$9276$new_n2194)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11126 (
        .A($abc$9276$new_n737), .B($abc$9276$new_n2194), .Y($abc$9276$new_n2195)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11127 (
        .A($abc$9276$new_n2195), .Y($abc$9276$new_n2196)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11128 (
        .A(CPU.ALU.CO), .B($abc$9276$new_n2178), .Y($abc$9276$new_n2197)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11129 (
        .A($abc$9276$new_n2197), .Y($abc$9276$new_n2198)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11130 (
        .A($abc$9276$new_n1438), .B($abc$9276$new_n1481), .Y($abc$9276$new_n2199)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11131 (
        .A($abc$9276$new_n1451), .B($abc$9276$new_n2199), .X($abc$9276$new_n2200)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11132 (
        .A($abc$9276$new_n1879), .B($abc$9276$new_n2200), .X($abc$9276$new_n2201)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11133 (
        .A(CPU.shift), .B(CPU.inc), .X($abc$9276$new_n2202)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11134 (
        .A(CPU.shift), .B($abc$9276$new_n377), .Y($abc$9276$new_n2203)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11135 (
        .A($abc$9276$new_n2202), .B($abc$9276$new_n2203), .Y($abc$9276$new_n2204)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11136 (
        .A(CPU.rotate), .B($abc$9276$new_n2204), .X($abc$9276$new_n2205)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11137 (
        .A($abc$9276$new_n2185), .B($abc$9276$new_n2205), .Y($abc$9276$new_n2206)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11138 (
        .A($abc$9276$new_n1478), .B($abc$9276$new_n2206), .Y($abc$9276$new_n2207)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11139 (
        .A($abc$9276$new_n1978), .B($abc$9276$new_n2207), .Y($abc$9276$new_n2208)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11140 (
        .A($abc$9276$new_n2201), .B($abc$9276$new_n2208), .X($abc$9276$new_n2209)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11141 (
        .A($abc$9276$new_n2198), .B($abc$9276$new_n2209), .X($abc$9276$new_n2210)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11142 (
        .A($abc$9276$new_n2196), .B($abc$9276$new_n2210), .X($abc$9276$new_n2211)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11143 (
        .A($abc$9276$new_n2184), .B($abc$9276$new_n2211), .X($abc$9276$new_n2212)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11144 (
        .A(CPU.shift_right), .B($abc$9276$new_n2180), .Y($abc$9276$new_n2213)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11145 (
        .A($abc$9276$new_n2181), .B($abc$9276$new_n2213), .Y($abc$9276$new_n2214)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11146 (
        .A($abc$9276$new_n2214), .Y($abc$9276$new_n2215)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11147 (
        .A($abc$9276$new_n2212), .B($abc$9276$new_n2215), .X($abc$9276$new_n2216)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11148 (
        .A($abc$9276$new_n390), .B($abc$9276$new_n398), .Y($abc$9276$new_n2217)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11149 (
        .A($abc$9276$new_n1476), .B($abc$9276$new_n2217), .X($abc$9276$new_n2218)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11150 (
        .A($abc$9276$new_n1504), .B($abc$9276$new_n2218), .X($abc$9276$new_n2219)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11151 (
        .A($abc$9276$new_n404), .B($abc$9276$new_n2009), .X($abc$9276$new_n2220)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11152 (
        .A($abc$9276$new_n440), .B($abc$9276$new_n2220), .X($abc$9276$new_n2221)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11153 (
        .A($abc$9276$new_n2219), .B($abc$9276$new_n2221), .X($abc$9276$new_n2222)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11154 (
        .A(CPU.load_only), .B($abc$9276$new_n736), .X($abc$9276$new_n2223)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11155 (
        .A($abc$9276$new_n2223), .Y($abc$9276$new_n2224)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11156 (
        .A($abc$9276$new_n2222), .B($abc$9276$new_n2224), .X($abc$9276$new_n2225)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11157 (
        .A($abc$9276$new_n2225), .Y($abc$9276$new_n2226)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11158 (
        .A($abc$9276$new_n1673), .B($abc$9276$new_n2226), .X($abc$9276$new_n2227)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11159 (
        .A($abc$9276$new_n1438), .B($abc$9276$new_n1453), .Y($abc$9276$new_n2228)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11160 (
        .A($abc$9276$new_n1451), .B($abc$9276$new_n2228), .X($abc$9276$new_n2229)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11161 (
        .A($abc$9276$new_n1449), .B($abc$9276$new_n2229), .X($abc$9276$new_n2230)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11162 (
        .A($abc$9276$new_n737), .B($abc$9276$new_n2179), .X($abc$9276$new_n2231)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11163 (
        .A($abc$9276$new_n1001), .B($abc$9276$new_n1477), .Y($abc$9276$new_n2232)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11164 (
        .A($abc$9276$new_n991), .B($abc$9276$new_n2232), .X($abc$9276$new_n2233)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11165 (
        .A($abc$9276$new_n2231), .B($abc$9276$new_n2233), .X($abc$9276$new_n2234)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11166 (
        .A($abc$9276$new_n2230), .B($abc$9276$new_n2234), .X($abc$9276$new_n2235)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11167 (
        .A($abc$9276$new_n2222), .B($abc$9276$new_n2235), .X($abc$9276$new_n2236)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11168 (
        .A($abc$9276$new_n2236), .Y($abc$9276$new_n2237)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11169 (
        .A(CPU.load_only), .B(oeb_0), .Y($abc$9276$new_n2238)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11170 (
        .A($abc$9276$new_n736), .B($abc$9276$new_n2238), .X($abc$9276$new_n2239)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11171 (
        .A($abc$9276$new_n2236), .B($abc$9276$new_n2239), .Y($abc$9276$new_n2240)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11172 (
        .A(CPU.ALU.N), .B($abc$9276$new_n2230), .Y($abc$9276$new_n2241)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11173 (
        .A(CPU.DIMUX), .B($abc$9276$new_n2232), .Y($abc$9276$new_n2242)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11174 (
        .A($abc$9276$new_n1308), .B($abc$9276$new_n2242), .Y($abc$9276$new_n2243)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11175 (
        .A($abc$9276$new_n2243), .Y($abc$9276$new_n2244)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11176 (
        .A($abc$9276$new_n2241), .B($abc$9276$new_n2244), .Y($abc$9276$new_n2245)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11177 (
        .A($abc$9276$new_n2240), .B($abc$9276$new_n2245), .X($abc$9276$new_n2246)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11178 (
        .A($abc$9276$new_n2246), .Y($abc$9276$new_n2247)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11179 (
        .A($abc$9276$new_n2227), .B($abc$9276$new_n2247), .Y($abc$9276$new_n2248)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11180 (
        .A(CPU.op), .B($abc$9276$new_n2180), .Y($abc$9276$new_n2249)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11181 (
        .A($abc$9276$new_n2249), .Y($abc$9276$new_n2250)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11182 (
        .A(CPU.op), .B($abc$9276$new_n2180), .Y($abc$9276$new_n2251)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11183 (
        .A($abc$9276$new_n2251), .Y($abc$9276$new_n2252)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11184 (
        .A($abc$9276$new_n392), .B($abc$9276$new_n1919), .X($abc$9276$new_n2253)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11185 (
        .A($abc$9276$new_n1886), .B($abc$9276$new_n2253), .X($abc$9276$new_n2254)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11186 (
        .A($abc$9276$new_n978), .B($abc$9276$new_n2254), .X($abc$9276$new_n2255)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11187 (
        .A($abc$9276$new_n351), .B($abc$9276$new_n1478), .X($abc$9276$new_n2256)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11188 (
        .A($abc$9276$new_n2231), .B($abc$9276$new_n2256), .X($abc$9276$new_n2257)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11189 (
        .A($abc$9276$new_n2257), .Y($abc$9276$new_n2258)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11190 (
        .A($abc$9276$new_n2255), .B($abc$9276$new_n2258), .X($abc$9276$new_n2259)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11191 (
        .A($abc$9276$new_n2252), .B($abc$9276$new_n2259), .X($abc$9276$new_n2260)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11192 (
        .A($abc$9276$new_n2250), .B($abc$9276$new_n2259), .X($abc$9276$new_n2261)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11193 (
        .A($abc$9276$new_n2250), .B($abc$9276$new_n2260), .X($abc$9276$new_n2262)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11194 (
        .A($abc$9276$new_n1450), .B($abc$9276$new_n1477), .Y($abc$9276$new_n2263)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11195 (
        .A($abc$9276$new_n1445), .B($abc$9276$new_n2263), .X($abc$9276$new_n2264)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11196 (
        .A($abc$9276$new_n2179), .B($abc$9276$new_n2228), .X($abc$9276$new_n2265)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11197 (
        .A($abc$9276$new_n2264), .B($abc$9276$new_n2265), .X($abc$9276$new_n2266)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11198 (
        .A($abc$9276$new_n2004), .B($abc$9276$new_n2220), .X($abc$9276$new_n2267)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11199 (
        .A($abc$9276$new_n2266), .B($abc$9276$new_n2267), .X($abc$9276$new_n2268)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11200 (
        .A($abc$9276$new_n2219), .B($abc$9276$new_n2268), .X($abc$9276$new_n2269)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11201 (
        .A($abc$9276$new_n2269), .Y($abc$9276$new_n2270)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11202 (
        .A(CPU.DIMUX), .B($abc$9276$new_n2270), .Y($abc$9276$new_n2271)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11203 (
        .A(CPU.PC), .B($abc$9276$new_n1002), .Y($abc$9276$new_n2272)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11204 (
        .A($abc$9276$new_n2271), .B($abc$9276$new_n2272), .Y($abc$9276$new_n2273)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11205 (
        .A($abc$9276$new_n2273), .Y($abc$9276$new_n2274)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11206 (
        .A($abc$9276$new_n2261), .B($abc$9276$new_n2274), .X($abc$9276$new_n2275)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11207 (
        .A($abc$9276$new_n2260), .B($abc$9276$new_n2273), .X($abc$9276$new_n2276)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11208 (
        .A($abc$9276$new_n2275), .B($abc$9276$new_n2276), .Y($abc$9276$new_n2277)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11209 (
        .A($abc$9276$new_n2262), .B($abc$9276$new_n2277), .Y($abc$9276$new_n2278)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11210 (
        .A($abc$9276$new_n2248), .B($abc$9276$new_n2275), .X($abc$9276$new_n2279)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11211 (
        .A($abc$9276$new_n2279), .Y($abc$9276$new_n2280)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11212 (
        .A($abc$9276$new_n2248), .B($abc$9276$new_n2278), .Y($abc$9276$new_n2281)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11213 (
        .A($abc$9276$new_n2215), .B($abc$9276$new_n2281), .Y($abc$9276$new_n2282)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11214 (
        .A($abc$9276$new_n2280), .B($abc$9276$new_n2282), .X($abc$9276$new_n2283)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11215 (
        .A($abc$9276$new_n2216), .B($abc$9276$new_n2283), .Y($abc$9276$new_n2284)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11216 (
        .A($abc$9276$new_n2182), .B($abc$9276$new_n2255), .X($abc$9276$new_n2285)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11217 (
        .A(CPU.op), .B($abc$9276$new_n2180), .Y($abc$9276$new_n2286)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11218 (
        .A($abc$9276$new_n2285), .B($abc$9276$new_n2286), .Y($abc$9276$new_n2287)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11219 (
        .A(CPU.backwards), .B($abc$9276$new_n978), .Y($abc$9276$new_n2288)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11220 (
        .A(CPU.op), .B($abc$9276$new_n2180), .Y($abc$9276$new_n2289)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11221 (
        .A($abc$9276$new_n2288), .B($abc$9276$new_n2289), .Y($abc$9276$new_n2290)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11222 (
        .A($abc$9276$new_n2254), .B($abc$9276$new_n2290), .X($abc$9276$new_n2291)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11223 (
        .A($abc$9276$new_n2291), .Y($abc$9276$new_n2292)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11224 (
        .A($abc$9276$new_n2285), .B($abc$9276$new_n2292), .Y($abc$9276$new_n2293)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11225 (
        .A($abc$9276$new_n2287), .B($abc$9276$new_n2291), .X($abc$9276$new_n2294)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11226 (
        .A($abc$9276$new_n2273), .B($abc$9276$new_n2294), .Y($abc$9276$new_n2295)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11227 (
        .A($abc$9276$new_n2287), .B($abc$9276$new_n2292), .X($abc$9276$new_n2296)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11228 (
        .A($abc$9276$new_n2274), .B($abc$9276$new_n2296), .Y($abc$9276$new_n2297)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11229 (
        .A($abc$9276$new_n2295), .B($abc$9276$new_n2297), .Y($abc$9276$new_n2298)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11230 (
        .A($abc$9276$new_n2284), .B($abc$9276$new_n2298), .Y($abc$9276$new_n2299)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11231 (
        .A($abc$9276$new_n2286), .B($abc$9276$new_n2293), .X($abc$9276$new_n2300)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11232 (
        .A($abc$9276$new_n2300), .Y($abc$9276$new_n2301)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11233 (
        .A($abc$9276$new_n2298), .B($abc$9276$new_n2300), .Y($abc$9276$new_n2302)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11234 (
        .A($abc$9276$new_n2302), .Y($abc$9276$new_n2303)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11235 (
        .A($abc$9276$new_n2299), .B($abc$9276$new_n2302), .Y($abc$9276$new_n2304)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11236 (
        .A($abc$9276$new_n359), .B($abc$9276$new_n2304), .X($abc$9276$new_n2305)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11237 (
        .A($abc$9276$new_n2177), .B($abc$9276$new_n2305), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9087)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11238 (
        .A(in_35), .B(CPU.ALU.N), .X($abc$9276$new_n2307)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11239 (
        .A($abc$9276$new_n606), .B($abc$9276$new_n2269), .X($abc$9276$new_n2308)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11240 (
        .A(CPU.PC), .B($abc$9276$new_n1002), .Y($abc$9276$new_n2309)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11241 (
        .A($abc$9276$new_n2308), .B($abc$9276$new_n2309), .Y($abc$9276$new_n2310)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11242 (
        .A($abc$9276$new_n2310), .Y($abc$9276$new_n2311)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11243 (
        .A($abc$9276$new_n2296), .B($abc$9276$new_n2310), .X($abc$9276$new_n2312)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11244 (
        .A($abc$9276$new_n2294), .B($abc$9276$new_n2311), .X($abc$9276$new_n2313)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11245 (
        .A($abc$9276$new_n2312), .B($abc$9276$new_n2313), .Y($abc$9276$new_n2314)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11246 (
        .A($abc$9276$new_n2301), .B($abc$9276$new_n2314), .X($abc$9276$new_n2315)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11247 (
        .A($abc$9276$new_n1647), .B($abc$9276$new_n2226), .X($abc$9276$new_n2316)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11248 (
        .A(CPU.ADD), .B($abc$9276$new_n2230), .Y($abc$9276$new_n2317)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11249 (
        .A(CPU.DIMUX), .B($abc$9276$new_n2232), .Y($abc$9276$new_n2318)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11250 (
        .A($abc$9276$new_n1288), .B($abc$9276$new_n2318), .Y($abc$9276$new_n2319)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11251 (
        .A($abc$9276$new_n2239), .B($abc$9276$new_n2317), .Y($abc$9276$new_n2320)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11252 (
        .A($abc$9276$new_n2237), .B($abc$9276$new_n2320), .X($abc$9276$new_n2321)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11253 (
        .A($abc$9276$new_n2319), .B($abc$9276$new_n2321), .X($abc$9276$new_n2322)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11254 (
        .A($abc$9276$new_n2322), .Y($abc$9276$new_n2323)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11255 (
        .A($abc$9276$new_n2316), .B($abc$9276$new_n2323), .Y($abc$9276$new_n2324)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11256 (
        .A($abc$9276$new_n2324), .Y($abc$9276$new_n2325)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11257 (
        .A($abc$9276$new_n2261), .B($abc$9276$new_n2311), .X($abc$9276$new_n2326)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11258 (
        .A($abc$9276$new_n2325), .B($abc$9276$new_n2326), .Y($abc$9276$new_n2327)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11259 (
        .A($abc$9276$new_n2327), .Y($abc$9276$new_n2328)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11260 (
        .A($abc$9276$new_n2260), .B($abc$9276$new_n2310), .X($abc$9276$new_n2329)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11261 (
        .A($abc$9276$new_n2326), .B($abc$9276$new_n2329), .Y($abc$9276$new_n2330)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11262 (
        .A($abc$9276$new_n2262), .B($abc$9276$new_n2330), .Y($abc$9276$new_n2331)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11263 (
        .A($abc$9276$new_n2325), .B($abc$9276$new_n2331), .X($abc$9276$new_n2332)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11264 (
        .A($abc$9276$new_n2214), .B($abc$9276$new_n2248), .Y($abc$9276$new_n2333)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11265 (
        .A($abc$9276$new_n2215), .B($abc$9276$new_n2332), .Y($abc$9276$new_n2334)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11266 (
        .A($abc$9276$new_n2328), .B($abc$9276$new_n2334), .X($abc$9276$new_n2335)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11267 (
        .A($abc$9276$new_n2333), .B($abc$9276$new_n2335), .Y($abc$9276$new_n2336)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11268 (
        .A($abc$9276$new_n2315), .B($abc$9276$new_n2336), .Y($abc$9276$new_n2337)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11269 (
        .A($abc$9276$new_n586), .B($abc$9276$new_n2269), .X($abc$9276$new_n2338)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11270 (
        .A(CPU.PC), .B($abc$9276$new_n1002), .Y($abc$9276$new_n2339)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11271 (
        .A($abc$9276$new_n2338), .B($abc$9276$new_n2339), .Y($abc$9276$new_n2340)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11272 (
        .A($abc$9276$new_n2340), .Y($abc$9276$new_n2341)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11273 (
        .A($abc$9276$new_n2294), .B($abc$9276$new_n2340), .Y($abc$9276$new_n2342)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11274 (
        .A($abc$9276$new_n2296), .B($abc$9276$new_n2341), .Y($abc$9276$new_n2343)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11275 (
        .A($abc$9276$new_n2342), .B($abc$9276$new_n2343), .Y($abc$9276$new_n2344)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11276 (
        .A($abc$9276$new_n2300), .B($abc$9276$new_n2344), .Y($abc$9276$new_n2345)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11277 (
        .A($abc$9276$new_n2345), .Y($abc$9276$new_n2346)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11278 (
        .A($abc$9276$new_n1621), .B($abc$9276$new_n2226), .X($abc$9276$new_n2347)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11279 (
        .A(CPU.ADD), .B($abc$9276$new_n2230), .Y($abc$9276$new_n2348)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11280 (
        .A(CPU.DIMUX), .B($abc$9276$new_n2232), .Y($abc$9276$new_n2349)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11281 (
        .A($abc$9276$new_n1270), .B($abc$9276$new_n2349), .Y($abc$9276$new_n2350)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11282 (
        .A($abc$9276$new_n2350), .Y($abc$9276$new_n2351)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11283 (
        .A($abc$9276$new_n2348), .B($abc$9276$new_n2351), .Y($abc$9276$new_n2352)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11284 (
        .A($abc$9276$new_n2240), .B($abc$9276$new_n2352), .X($abc$9276$new_n2353)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11285 (
        .A($abc$9276$new_n2353), .Y($abc$9276$new_n2354)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11286 (
        .A($abc$9276$new_n2347), .B($abc$9276$new_n2354), .Y($abc$9276$new_n2355)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11287 (
        .A($abc$9276$new_n2261), .B($abc$9276$new_n2341), .X($abc$9276$new_n2356)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11288 (
        .A($abc$9276$new_n2260), .B($abc$9276$new_n2340), .X($abc$9276$new_n2357)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11289 (
        .A($abc$9276$new_n2356), .B($abc$9276$new_n2357), .Y($abc$9276$new_n2358)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11290 (
        .A($abc$9276$new_n2262), .B($abc$9276$new_n2358), .Y($abc$9276$new_n2359)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11291 (
        .A($abc$9276$new_n2355), .B($abc$9276$new_n2356), .X($abc$9276$new_n2360)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11292 (
        .A($abc$9276$new_n2355), .B($abc$9276$new_n2359), .Y($abc$9276$new_n2361)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11293 (
        .A($abc$9276$new_n2360), .B($abc$9276$new_n2361), .Y($abc$9276$new_n2362)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11294 (
        .A($abc$9276$new_n2214), .B($abc$9276$new_n2362), .X($abc$9276$new_n2363)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11295 (
        .A($abc$9276$new_n2215), .B($abc$9276$new_n2324), .X($abc$9276$new_n2364)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11296 (
        .A($abc$9276$new_n2363), .B($abc$9276$new_n2364), .Y($abc$9276$new_n2365)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11297 (
        .A($abc$9276$new_n2346), .B($abc$9276$new_n2365), .X($abc$9276$new_n2366)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11298 (
        .A(CPU.DIMUX), .B($abc$9276$new_n2270), .Y($abc$9276$new_n2367)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11299 (
        .A(CPU.PC), .B($abc$9276$new_n1002), .Y($abc$9276$new_n2368)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11300 (
        .A($abc$9276$new_n2367), .B($abc$9276$new_n2368), .Y($abc$9276$new_n2369)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11301 (
        .A($abc$9276$new_n2369), .Y($abc$9276$new_n2370)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11302 (
        .A($abc$9276$new_n2296), .B($abc$9276$new_n2369), .X($abc$9276$new_n2371)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11303 (
        .A($abc$9276$new_n2294), .B($abc$9276$new_n2370), .X($abc$9276$new_n2372)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11304 (
        .A($abc$9276$new_n2371), .B($abc$9276$new_n2372), .Y($abc$9276$new_n2373)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11305 (
        .A($abc$9276$new_n2301), .B($abc$9276$new_n2373), .X($abc$9276$new_n2374)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11306 (
        .A($abc$9276$new_n1595), .B($abc$9276$new_n2226), .X($abc$9276$new_n2375)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11307 (
        .A(CPU.ADD), .B($abc$9276$new_n2230), .Y($abc$9276$new_n2376)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11308 (
        .A(CPU.DIMUX), .B($abc$9276$new_n2232), .Y($abc$9276$new_n2377)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11309 (
        .A($abc$9276$new_n1251), .B($abc$9276$new_n2377), .Y($abc$9276$new_n2378)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11310 (
        .A($abc$9276$new_n2378), .Y($abc$9276$new_n2379)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11311 (
        .A($abc$9276$new_n2376), .B($abc$9276$new_n2379), .Y($abc$9276$new_n2380)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11312 (
        .A($abc$9276$new_n2240), .B($abc$9276$new_n2380), .X($abc$9276$new_n2381)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11313 (
        .A($abc$9276$new_n2381), .Y($abc$9276$new_n2382)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11314 (
        .A($abc$9276$new_n2375), .B($abc$9276$new_n2382), .Y($abc$9276$new_n2383)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11315 (
        .A($abc$9276$new_n2261), .B($abc$9276$new_n2370), .X($abc$9276$new_n2384)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11316 (
        .A($abc$9276$new_n2384), .Y($abc$9276$new_n2385)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11317 (
        .A($abc$9276$new_n2260), .B($abc$9276$new_n2369), .X($abc$9276$new_n2386)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11318 (
        .A($abc$9276$new_n2384), .B($abc$9276$new_n2386), .Y($abc$9276$new_n2387)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11319 (
        .A($abc$9276$new_n2262), .B($abc$9276$new_n2387), .Y($abc$9276$new_n2388)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11320 (
        .A($abc$9276$new_n2388), .Y($abc$9276$new_n2389)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11321 (
        .A($abc$9276$new_n2383), .B($abc$9276$new_n2389), .Y($abc$9276$new_n2390)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11322 (
        .A($abc$9276$new_n2383), .B($abc$9276$new_n2385), .X($abc$9276$new_n2391)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11323 (
        .A($abc$9276$new_n2391), .Y($abc$9276$new_n2392)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11324 (
        .A($abc$9276$new_n2214), .B($abc$9276$new_n2355), .Y($abc$9276$new_n2393)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11325 (
        .A($abc$9276$new_n2215), .B($abc$9276$new_n2390), .Y($abc$9276$new_n2394)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11326 (
        .A($abc$9276$new_n2392), .B($abc$9276$new_n2394), .X($abc$9276$new_n2395)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11327 (
        .A($abc$9276$new_n2393), .B($abc$9276$new_n2395), .Y($abc$9276$new_n2396)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11328 (
        .A($abc$9276$new_n2374), .B($abc$9276$new_n2396), .Y($abc$9276$new_n2397)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11329 (
        .A($abc$9276$new_n545), .B($abc$9276$new_n2269), .X($abc$9276$new_n2398)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11330 (
        .A(CPU.PC), .B($abc$9276$new_n1002), .Y($abc$9276$new_n2399)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11331 (
        .A($abc$9276$new_n2398), .B($abc$9276$new_n2399), .Y($abc$9276$new_n2400)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11332 (
        .A($abc$9276$new_n2400), .Y($abc$9276$new_n2401)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11333 (
        .A($abc$9276$new_n2294), .B($abc$9276$new_n2400), .Y($abc$9276$new_n2402)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11334 (
        .A($abc$9276$new_n2296), .B($abc$9276$new_n2401), .Y($abc$9276$new_n2403)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11335 (
        .A($abc$9276$new_n2402), .B($abc$9276$new_n2403), .Y($abc$9276$new_n2404)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11336 (
        .A($abc$9276$new_n2300), .B($abc$9276$new_n2404), .Y($abc$9276$new_n2405)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11337 (
        .A($abc$9276$new_n2405), .Y($abc$9276$new_n2406)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11338 (
        .A($abc$9276$new_n1569), .B($abc$9276$new_n2226), .X($abc$9276$new_n2407)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11339 (
        .A(CPU.ADD), .B($abc$9276$new_n2230), .Y($abc$9276$new_n2408)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11340 (
        .A(CPU.DIMUX), .B($abc$9276$new_n2232), .Y($abc$9276$new_n2409)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11341 (
        .A($abc$9276$new_n1230), .B($abc$9276$new_n2409), .Y($abc$9276$new_n2410)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11342 (
        .A($abc$9276$new_n2410), .Y($abc$9276$new_n2411)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11343 (
        .A($abc$9276$new_n2408), .B($abc$9276$new_n2411), .Y($abc$9276$new_n2412)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11344 (
        .A($abc$9276$new_n2240), .B($abc$9276$new_n2412), .X($abc$9276$new_n2413)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11345 (
        .A($abc$9276$new_n2413), .Y($abc$9276$new_n2414)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11346 (
        .A($abc$9276$new_n2407), .B($abc$9276$new_n2414), .Y($abc$9276$new_n2415)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11347 (
        .A($abc$9276$new_n2261), .B($abc$9276$new_n2401), .X($abc$9276$new_n2416)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11348 (
        .A($abc$9276$new_n2260), .B($abc$9276$new_n2400), .X($abc$9276$new_n2417)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11349 (
        .A($abc$9276$new_n2416), .B($abc$9276$new_n2417), .Y($abc$9276$new_n2418)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11350 (
        .A($abc$9276$new_n2262), .B($abc$9276$new_n2418), .Y($abc$9276$new_n2419)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11351 (
        .A($abc$9276$new_n2415), .B($abc$9276$new_n2416), .X($abc$9276$new_n2420)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11352 (
        .A($abc$9276$new_n2415), .B($abc$9276$new_n2419), .Y($abc$9276$new_n2421)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11353 (
        .A($abc$9276$new_n2420), .B($abc$9276$new_n2421), .Y($abc$9276$new_n2422)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11354 (
        .A($abc$9276$new_n2214), .B($abc$9276$new_n2422), .X($abc$9276$new_n2423)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11355 (
        .A($abc$9276$new_n2215), .B($abc$9276$new_n2383), .X($abc$9276$new_n2424)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11356 (
        .A($abc$9276$new_n2423), .B($abc$9276$new_n2424), .Y($abc$9276$new_n2425)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11357 (
        .A($abc$9276$new_n2406), .B($abc$9276$new_n2425), .X($abc$9276$new_n2426)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11358 (
        .A($abc$9276$new_n2404), .B($abc$9276$new_n2425), .Y($abc$9276$new_n2427)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11359 (
        .A($abc$9276$new_n2426), .B($abc$9276$new_n2427), .Y($abc$9276$new_n2428)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11360 (
        .A($abc$9276$new_n2428), .Y($abc$9276$new_n2429)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11361 (
        .A($abc$9276$new_n525), .B($abc$9276$new_n2269), .X($abc$9276$new_n2430)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11362 (
        .A(CPU.PC), .B($abc$9276$new_n1002), .Y($abc$9276$new_n2431)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11363 (
        .A($abc$9276$new_n2430), .B($abc$9276$new_n2431), .Y($abc$9276$new_n2432)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11364 (
        .A($abc$9276$new_n2432), .Y($abc$9276$new_n2433)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11365 (
        .A($abc$9276$new_n2294), .B($abc$9276$new_n2432), .Y($abc$9276$new_n2434)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11366 (
        .A($abc$9276$new_n2296), .B($abc$9276$new_n2433), .Y($abc$9276$new_n2435)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11367 (
        .A($abc$9276$new_n2434), .B($abc$9276$new_n2435), .Y($abc$9276$new_n2436)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11368 (
        .A($abc$9276$new_n2300), .B($abc$9276$new_n2436), .Y($abc$9276$new_n2437)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11369 (
        .A($abc$9276$new_n2437), .Y($abc$9276$new_n2438)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11370 (
        .A($abc$9276$new_n1544), .B($abc$9276$new_n2226), .X($abc$9276$new_n2439)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11371 (
        .A(CPU.ADD), .B($abc$9276$new_n2230), .Y($abc$9276$new_n2440)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11372 (
        .A(CPU.DIMUX), .B($abc$9276$new_n2232), .Y($abc$9276$new_n2441)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11373 (
        .A($abc$9276$new_n2239), .B($abc$9276$new_n2441), .Y($abc$9276$new_n2442)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11374 (
        .A($abc$9276$new_n1211), .B($abc$9276$new_n2442), .X($abc$9276$new_n2443)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11375 (
        .A($abc$9276$new_n2443), .Y($abc$9276$new_n2444)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11376 (
        .A($abc$9276$new_n2440), .B($abc$9276$new_n2444), .Y($abc$9276$new_n2445)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11377 (
        .A($abc$9276$new_n2237), .B($abc$9276$new_n2445), .X($abc$9276$new_n2446)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11378 (
        .A($abc$9276$new_n2446), .Y($abc$9276$new_n2447)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11379 (
        .A($abc$9276$new_n2439), .B($abc$9276$new_n2447), .Y($abc$9276$new_n2448)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11380 (
        .A($abc$9276$new_n2261), .B($abc$9276$new_n2433), .X($abc$9276$new_n2449)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11381 (
        .A($abc$9276$new_n2260), .B($abc$9276$new_n2432), .X($abc$9276$new_n2450)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11382 (
        .A($abc$9276$new_n2449), .B($abc$9276$new_n2450), .Y($abc$9276$new_n2451)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11383 (
        .A($abc$9276$new_n2262), .B($abc$9276$new_n2451), .Y($abc$9276$new_n2452)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11384 (
        .A($abc$9276$new_n2448), .B($abc$9276$new_n2449), .X($abc$9276$new_n2453)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11385 (
        .A($abc$9276$new_n2448), .B($abc$9276$new_n2452), .Y($abc$9276$new_n2454)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11386 (
        .A($abc$9276$new_n2453), .B($abc$9276$new_n2454), .Y($abc$9276$new_n2455)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11387 (
        .A($abc$9276$new_n2214), .B($abc$9276$new_n2455), .X($abc$9276$new_n2456)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11388 (
        .A($abc$9276$new_n2215), .B($abc$9276$new_n2415), .X($abc$9276$new_n2457)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11389 (
        .A($abc$9276$new_n2456), .B($abc$9276$new_n2457), .Y($abc$9276$new_n2458)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11390 (
        .A($abc$9276$new_n2438), .B($abc$9276$new_n2458), .X($abc$9276$new_n2459)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11391 (
        .A($abc$9276$new_n505), .B($abc$9276$new_n2269), .X($abc$9276$new_n2460)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11392 (
        .A(CPU.PC), .B($abc$9276$new_n1002), .Y($abc$9276$new_n2461)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11393 (
        .A($abc$9276$new_n2460), .B($abc$9276$new_n2461), .Y($abc$9276$new_n2462)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11394 (
        .A($abc$9276$new_n2462), .Y($abc$9276$new_n2463)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11395 (
        .A($abc$9276$new_n2296), .B($abc$9276$new_n2462), .X($abc$9276$new_n2464)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11396 (
        .A($abc$9276$new_n2294), .B($abc$9276$new_n2463), .X($abc$9276$new_n2465)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11397 (
        .A($abc$9276$new_n2464), .B($abc$9276$new_n2465), .Y($abc$9276$new_n2466)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11398 (
        .A($abc$9276$new_n2301), .B($abc$9276$new_n2466), .X($abc$9276$new_n2467)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11399 (
        .A($abc$9276$new_n1521), .B($abc$9276$new_n2226), .X($abc$9276$new_n2468)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11400 (
        .A(CPU.ADD), .B($abc$9276$new_n2230), .Y($abc$9276$new_n2469)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11401 (
        .A(CPU.DIMUX), .B($abc$9276$new_n2232), .Y($abc$9276$new_n2470)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11402 (
        .A($abc$9276$new_n1190), .B($abc$9276$new_n2236), .Y($abc$9276$new_n2471)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11403 (
        .A($abc$9276$new_n2239), .B($abc$9276$new_n2470), .Y($abc$9276$new_n2472)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11404 (
        .A($abc$9276$new_n2472), .Y($abc$9276$new_n2473)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11405 (
        .A($abc$9276$new_n2469), .B($abc$9276$new_n2473), .Y($abc$9276$new_n2474)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11406 (
        .A($abc$9276$new_n2471), .B($abc$9276$new_n2474), .X($abc$9276$new_n2475)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11407 (
        .A($abc$9276$new_n2475), .Y($abc$9276$new_n2476)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11408 (
        .A($abc$9276$new_n2468), .B($abc$9276$new_n2476), .Y($abc$9276$new_n2477)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11409 (
        .A($abc$9276$new_n2261), .B($abc$9276$new_n2463), .X($abc$9276$new_n2478)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11410 (
        .A($abc$9276$new_n2260), .B($abc$9276$new_n2462), .X($abc$9276$new_n2479)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11411 (
        .A($abc$9276$new_n2478), .B($abc$9276$new_n2479), .Y($abc$9276$new_n2480)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11412 (
        .A($abc$9276$new_n2262), .B($abc$9276$new_n2480), .Y($abc$9276$new_n2481)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11413 (
        .A($abc$9276$new_n2477), .B($abc$9276$new_n2481), .Y($abc$9276$new_n2482)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11414 (
        .A($abc$9276$new_n2477), .B($abc$9276$new_n2478), .X($abc$9276$new_n2483)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11415 (
        .A($abc$9276$new_n2482), .B($abc$9276$new_n2483), .Y($abc$9276$new_n2484)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11416 (
        .A($abc$9276$new_n2215), .B($abc$9276$new_n2484), .Y($abc$9276$new_n2485)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11417 (
        .A($abc$9276$new_n2214), .B($abc$9276$new_n2448), .Y($abc$9276$new_n2486)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11418 (
        .A($abc$9276$new_n2485), .B($abc$9276$new_n2486), .Y($abc$9276$new_n2487)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11419 (
        .A($abc$9276$new_n2467), .B($abc$9276$new_n2487), .Y($abc$9276$new_n2488)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11420 (
        .A($abc$9276$new_n487), .B($abc$9276$new_n2269), .X($abc$9276$new_n2489)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11421 (
        .A(CPU.PC), .B($abc$9276$new_n1002), .Y($abc$9276$new_n2490)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11422 (
        .A($abc$9276$new_n2489), .B($abc$9276$new_n2490), .Y($abc$9276$new_n2491)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11423 (
        .A($abc$9276$new_n2491), .Y($abc$9276$new_n2492)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11424 (
        .A($abc$9276$new_n2296), .B($abc$9276$new_n2491), .X($abc$9276$new_n2493)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11425 (
        .A($abc$9276$new_n2294), .B($abc$9276$new_n2492), .X($abc$9276$new_n2494)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11426 (
        .A($abc$9276$new_n2493), .B($abc$9276$new_n2494), .Y($abc$9276$new_n2495)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11427 (
        .A($abc$9276$new_n2301), .B($abc$9276$new_n2495), .X($abc$9276$new_n2496)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11428 (
        .A($abc$9276$new_n2214), .B($abc$9276$new_n2477), .Y($abc$9276$new_n2497)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11429 (
        .A($abc$9276$new_n1436), .B($abc$9276$new_n2225), .Y($abc$9276$new_n2498)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11430 (
        .A(CPU.ADD), .B($abc$9276$new_n2230), .Y($abc$9276$new_n2499)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11431 (
        .A(CPU.DIMUX), .B($abc$9276$new_n2232), .Y($abc$9276$new_n2500)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11432 (
        .A($abc$9276$new_n1170), .B($abc$9276$new_n2500), .Y($abc$9276$new_n2501)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11433 (
        .A($abc$9276$new_n2501), .Y($abc$9276$new_n2502)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11434 (
        .A($abc$9276$new_n2499), .B($abc$9276$new_n2502), .Y($abc$9276$new_n2503)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11435 (
        .A($abc$9276$new_n2240), .B($abc$9276$new_n2503), .X($abc$9276$new_n2504)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11436 (
        .A($abc$9276$new_n2504), .Y($abc$9276$new_n2505)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11437 (
        .A($abc$9276$new_n2498), .B($abc$9276$new_n2505), .Y($abc$9276$new_n2506)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11438 (
        .A($abc$9276$new_n2261), .B($abc$9276$new_n2492), .X($abc$9276$new_n2507)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11439 (
        .A($abc$9276$new_n2260), .B($abc$9276$new_n2491), .X($abc$9276$new_n2508)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11440 (
        .A($abc$9276$new_n2507), .B($abc$9276$new_n2508), .Y($abc$9276$new_n2509)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11441 (
        .A($abc$9276$new_n2262), .B($abc$9276$new_n2509), .Y($abc$9276$new_n2510)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11442 (
        .A($abc$9276$new_n2506), .B($abc$9276$new_n2507), .X($abc$9276$new_n2511)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11443 (
        .A($abc$9276$new_n2506), .B($abc$9276$new_n2510), .Y($abc$9276$new_n2512)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11444 (
        .A($abc$9276$new_n2511), .B($abc$9276$new_n2512), .Y($abc$9276$new_n2513)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11445 (
        .A($abc$9276$new_n2215), .B($abc$9276$new_n2513), .Y($abc$9276$new_n2514)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11446 (
        .A($abc$9276$new_n2497), .B($abc$9276$new_n2514), .Y($abc$9276$new_n2515)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11447 (
        .A($abc$9276$new_n2496), .B($abc$9276$new_n2515), .Y($abc$9276$new_n2516)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11448 (
        .A($abc$9276$new_n2495), .B($abc$9276$new_n2515), .X($abc$9276$new_n2517)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11449 (
        .A($abc$9276$new_n2516), .B($abc$9276$new_n2517), .Y($abc$9276$new_n2518)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11450 (
        .A($abc$9276$new_n2287), .B($abc$9276$new_n2293), .Y($abc$9276$new_n2519)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11451 (
        .A($abc$9276$new_n2215), .B($abc$9276$new_n2519), .Y($abc$9276$new_n2520)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11452 (
        .A($abc$9276$new_n2212), .B($abc$9276$new_n2520), .X($abc$9276$new_n2521)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11453 (
        .A($abc$9276$new_n377), .B($abc$9276$new_n2520), .Y($abc$9276$new_n2522)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11454 (
        .A($abc$9276$new_n2521), .B($abc$9276$new_n2522), .Y($abc$9276$new_n2523)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11455 (
        .A($abc$9276$new_n2518), .B($abc$9276$new_n2523), .X($abc$9276$new_n2524)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11456 (
        .A($abc$9276$new_n2516), .B($abc$9276$new_n2524), .Y($abc$9276$new_n2525)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11457 (
        .A($abc$9276$new_n2466), .B($abc$9276$new_n2487), .X($abc$9276$new_n2526)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11458 (
        .A($abc$9276$new_n2488), .B($abc$9276$new_n2526), .Y($abc$9276$new_n2527)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11459 (
        .A($abc$9276$new_n2527), .Y($abc$9276$new_n2528)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11460 (
        .A($abc$9276$new_n2525), .B($abc$9276$new_n2528), .Y($abc$9276$new_n2529)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11461 (
        .A($abc$9276$new_n2488), .B($abc$9276$new_n2529), .Y($abc$9276$new_n2530)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11462 (
        .A($abc$9276$new_n2436), .B($abc$9276$new_n2458), .Y($abc$9276$new_n2531)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11463 (
        .A($abc$9276$new_n2459), .B($abc$9276$new_n2531), .Y($abc$9276$new_n2532)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11464 (
        .A($abc$9276$new_n2532), .Y($abc$9276$new_n2533)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11465 (
        .A($abc$9276$new_n2530), .B($abc$9276$new_n2533), .Y($abc$9276$new_n2534)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11466 (
        .A($abc$9276$new_n2459), .B($abc$9276$new_n2534), .Y($abc$9276$new_n2535)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11467 (
        .A($abc$9276$new_n2429), .B($abc$9276$new_n2535), .Y($abc$9276$new_n2536)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11468 (
        .A($abc$9276$new_n2429), .B($abc$9276$new_n2535), .X($abc$9276$new_n2537)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11469 (
        .A($abc$9276$new_n2536), .B($abc$9276$new_n2537), .Y($abc$9276$new_n2538)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11470 (
        .A(CPU.adc_bcd), .B($abc$9276$new_n737), .Y($abc$9276$new_n2539)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11471 (
        .A($abc$9276$new_n2539), .Y($abc$9276$new_n2540)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11472 (
        .A($abc$9276$new_n2530), .B($abc$9276$new_n2533), .X($abc$9276$new_n2541)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11473 (
        .A($abc$9276$new_n2534), .B($abc$9276$new_n2541), .Y($abc$9276$new_n2542)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11474 (
        .A($abc$9276$new_n2525), .B($abc$9276$new_n2528), .X($abc$9276$new_n2543)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11475 (
        .A($abc$9276$new_n2529), .B($abc$9276$new_n2543), .Y($abc$9276$new_n2544)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11476 (
        .A($abc$9276$new_n2542), .B($abc$9276$new_n2544), .Y($abc$9276$new_n2545)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11477 (
        .A($abc$9276$new_n2540), .B($abc$9276$new_n2545), .Y($abc$9276$new_n2546)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11478 (
        .A($abc$9276$new_n2538), .B($abc$9276$new_n2546), .X($abc$9276$new_n2547)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11479 (
        .A($abc$9276$new_n2426), .B($abc$9276$new_n2536), .Y($abc$9276$new_n2548)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11480 (
        .A($abc$9276$new_n2548), .Y($abc$9276$new_n2549)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11481 (
        .A($abc$9276$new_n2547), .B($abc$9276$new_n2549), .Y($abc$9276$new_n2550)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11482 (
        .A($abc$9276$new_n2373), .B($abc$9276$new_n2396), .X($abc$9276$new_n2551)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11483 (
        .A($abc$9276$new_n2397), .B($abc$9276$new_n2551), .Y($abc$9276$new_n2552)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11484 (
        .A($abc$9276$new_n2552), .Y($abc$9276$new_n2553)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11485 (
        .A($abc$9276$new_n2550), .B($abc$9276$new_n2553), .Y($abc$9276$new_n2554)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11486 (
        .A($abc$9276$new_n2397), .B($abc$9276$new_n2554), .Y($abc$9276$new_n2555)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11487 (
        .A($abc$9276$new_n2344), .B($abc$9276$new_n2365), .Y($abc$9276$new_n2556)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11488 (
        .A($abc$9276$new_n2366), .B($abc$9276$new_n2556), .Y($abc$9276$new_n2557)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11489 (
        .A($abc$9276$new_n2557), .Y($abc$9276$new_n2558)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11490 (
        .A($abc$9276$new_n2555), .B($abc$9276$new_n2558), .Y($abc$9276$new_n2559)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11491 (
        .A($abc$9276$new_n2366), .B($abc$9276$new_n2559), .Y($abc$9276$new_n2560)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11492 (
        .A($abc$9276$new_n2314), .B($abc$9276$new_n2336), .X($abc$9276$new_n2561)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11493 (
        .A($abc$9276$new_n2337), .B($abc$9276$new_n2561), .Y($abc$9276$new_n2562)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11494 (
        .A($abc$9276$new_n2562), .Y($abc$9276$new_n2563)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11495 (
        .A($abc$9276$new_n2560), .B($abc$9276$new_n2563), .Y($abc$9276$new_n2564)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11496 (
        .A($abc$9276$new_n2337), .B($abc$9276$new_n2564), .Y($abc$9276$new_n2565)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11497 (
        .A($abc$9276$new_n2284), .B($abc$9276$new_n2303), .X($abc$9276$new_n2566)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11498 (
        .A($abc$9276$new_n2566), .Y($abc$9276$new_n2567)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11499 (
        .A($abc$9276$new_n2299), .B($abc$9276$new_n2566), .Y($abc$9276$new_n2568)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11500 (
        .A($abc$9276$new_n2565), .B($abc$9276$new_n2568), .Y($abc$9276$new_n2569)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11501 (
        .A($abc$9276$new_n2565), .B($abc$9276$new_n2568), .X($abc$9276$new_n2570)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11502 (
        .A($abc$9276$new_n2569), .B($abc$9276$new_n2570), .Y($abc$9276$new_n2571)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11503 (
        .A($abc$9276$new_n359), .B($abc$9276$new_n2571), .X($abc$9276$new_n2572)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11504 (
        .A($abc$9276$new_n2307), .B($abc$9276$new_n2572), .Y($abc$9276$new_n2573)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11505 (
        .A($abc$9276$new_n2573), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9089)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11506 (
        .A($abc$9276$new_n359), .B(CPU.ALU.HC), .Y($abc$9276$new_n2575)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11507 (
        .A(in_35), .B($abc$9276$new_n2550), .Y($abc$9276$new_n2576)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11508 (
        .A($abc$9276$new_n2575), .B($abc$9276$new_n2576), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9091)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11509 (
        .A($abc$9276$new_n2518), .B($abc$9276$new_n2523), .Y($abc$9276$new_n2578)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11510 (
        .A($abc$9276$new_n2524), .B($abc$9276$new_n2578), .Y($abc$9276$new_n2579)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11511 (
        .A(in_35), .B($abc$9276$new_n2579), .Y($abc$9276$new_n2580)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11512 (
        .A(in_35), .B(CPU.ADD), .X($abc$9276$new_n2581)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11513 (
        .A($abc$9276$new_n2580), .B($abc$9276$new_n2581), .Y($abc$9276$new_n2582)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11514 (
        .A($abc$9276$new_n2582), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9093)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11515 (
        .A(in_35), .B(CPU.ADD), .X($abc$9276$new_n2584)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11516 (
        .A(in_35), .B($abc$9276$new_n2544), .Y($abc$9276$new_n2585)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11517 (
        .A($abc$9276$new_n2584), .B($abc$9276$new_n2585), .Y($abc$9276$new_n2586)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11518 (
        .A($abc$9276$new_n2586), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9095)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11519 (
        .A(in_35), .B(CPU.ADD), .X($abc$9276$new_n2588)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11520 (
        .A(in_35), .B($abc$9276$new_n2542), .Y($abc$9276$new_n2589)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11521 (
        .A($abc$9276$new_n2588), .B($abc$9276$new_n2589), .Y($abc$9276$new_n2590)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11522 (
        .A($abc$9276$new_n2590), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9097)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11523 (
        .A(in_35), .B(CPU.ADD), .X($abc$9276$new_n2592)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11524 (
        .A(in_35), .B($abc$9276$new_n2538), .Y($abc$9276$new_n2593)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11525 (
        .A($abc$9276$new_n2592), .B($abc$9276$new_n2593), .Y($abc$9276$new_n2594)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11526 (
        .A($abc$9276$new_n2594), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9099)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11527 (
        .A($abc$9276$new_n2550), .B($abc$9276$new_n2553), .X($abc$9276$new_n2596)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11528 (
        .A($abc$9276$new_n2554), .B($abc$9276$new_n2596), .Y($abc$9276$new_n2597)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11529 (
        .A(in_35), .B($abc$9276$new_n2597), .Y($abc$9276$new_n2598)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11530 (
        .A(in_35), .B(CPU.ADD), .X($abc$9276$new_n2599)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11531 (
        .A($abc$9276$new_n2598), .B($abc$9276$new_n2599), .Y($abc$9276$new_n2600)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11532 (
        .A($abc$9276$new_n2600), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9101)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11533 (
        .A($abc$9276$new_n2555), .B($abc$9276$new_n2558), .X($abc$9276$new_n2602)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11534 (
        .A($abc$9276$new_n2559), .B($abc$9276$new_n2602), .Y($abc$9276$new_n2603)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11535 (
        .A(in_35), .B(CPU.ADD), .X($abc$9276$new_n2604)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11536 (
        .A(in_35), .B($abc$9276$new_n2603), .Y($abc$9276$new_n2605)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11537 (
        .A($abc$9276$new_n2604), .B($abc$9276$new_n2605), .Y($abc$9276$new_n2606)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11538 (
        .A($abc$9276$new_n2606), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9103)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11539 (
        .A($abc$9276$new_n2560), .B($abc$9276$new_n2563), .X($abc$9276$new_n2608)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11540 (
        .A($abc$9276$new_n2564), .B($abc$9276$new_n2608), .Y($abc$9276$new_n2609)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11541 (
        .A(in_35), .B(CPU.ADD), .X($abc$9276$new_n2610)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11542 (
        .A(in_35), .B($abc$9276$new_n2609), .Y($abc$9276$new_n2611)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11543 (
        .A($abc$9276$new_n2610), .B($abc$9276$new_n2611), .Y($abc$9276$new_n2612)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11544 (
        .A($abc$9276$new_n2612), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9105)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11545 (
        .A($abc$9276$new_n359), .B(CPU.ALU.AI7), .Y($abc$9276$new_n2614)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11546 (
        .A(in_35), .B($abc$9276$new_n2248), .Y($abc$9276$new_n2615)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11547 (
        .A($abc$9276$new_n2614), .B($abc$9276$new_n2615), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9107)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11548 (
        .A(in_35), .B(CPU.ALU.CO), .X($abc$9276$new_n2617)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11549 (
        .A($abc$9276$new_n2215), .B($abc$9276$new_n2506), .X($abc$9276$new_n2618)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11550 (
        .A($abc$9276$new_n377), .B($abc$9276$new_n2213), .Y($abc$9276$new_n2619)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11551 (
        .A($abc$9276$new_n2618), .B($abc$9276$new_n2619), .Y($abc$9276$new_n2620)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11552 (
        .A($abc$9276$new_n2565), .B($abc$9276$new_n2567), .X($abc$9276$new_n2621)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11553 (
        .A($abc$9276$new_n2299), .B($abc$9276$new_n2621), .Y($abc$9276$new_n2622)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11554 (
        .A($abc$9276$new_n2620), .B($abc$9276$new_n2622), .X($abc$9276$new_n2623)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11555 (
        .A($abc$9276$new_n2620), .B($abc$9276$new_n2622), .Y($abc$9276$new_n2624)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11556 (
        .A($abc$9276$new_n2623), .B($abc$9276$new_n2624), .Y($abc$9276$new_n2625)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11557 (
        .A($abc$9276$new_n2603), .B($abc$9276$new_n2609), .Y($abc$9276$new_n2626)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11558 (
        .A($abc$9276$new_n2540), .B($abc$9276$new_n2626), .Y($abc$9276$new_n2627)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11559 (
        .A(in_35), .B($abc$9276$new_n2627), .Y($abc$9276$new_n2628)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11560 (
        .A($abc$9276$new_n2572), .B($abc$9276$new_n2628), .Y($abc$9276$new_n2629)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11561 (
        .A($abc$9276$new_n2625), .B($abc$9276$new_n2629), .Y($abc$9276$new_n2630)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11562 (
        .A($abc$9276$new_n2617), .B($abc$9276$new_n2630), .Y($abc$9276$new_n2631)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11563 (
        .A($abc$9276$new_n2631), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$9109)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11564 (
        .A($abc$9276$new_n350), .B($abc$9276$new_n410), .X($abc$9276$new_n2633)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11565 (
        .A(in_34), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9228), .Y($abc$9276$new_n2634)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11566 (
        .A($abc$9276$new_n351), .B($abc$9276$new_n2634), .X($abc$9276$new_n2635)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11567 (
        .A(CPU.NMI_edge), .B($abc$9276$new_n2634), .Y($abc$9276$new_n2636)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11568 (
        .A($abc$9276$new_n2635), .B($abc$9276$new_n2636), .Y($abc$9276$new_n2637)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11569 (
        .A($abc$9276$new_n2633), .B($abc$9276$new_n2637), .Y($abc$9276$new_n2638)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11570 (
        .A($abc$9276$new_n2638), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8887)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11571 (
        .A($abc$9276$new_n377), .B($abc$9276$new_n428), .X($abc$9276$new_n2640)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11572 (
        .A($abc$9276$new_n2640), .Y($abc$9276$new_n2641)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11573 (
        .A(CPU.res), .B($abc$9276$new_n428), .Y($abc$9276$new_n2642)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11574 (
        .A(rst_n), .B($abc$9276$new_n2642), .Y($abc$9276$new_n2643)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11575 (
        .A($abc$9276$new_n2641), .B($abc$9276$new_n2643), .X($abc$9276$auto$rtlil.cc:3205:MuxGate$8969)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11576 (
        .A($abc$9276$new_n752), .B($abc$9276$new_n1789), .Y($abc$9276$new_n2645)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11577 (
        .A(CPU.IRHOLD_valid), .B($abc$9276$new_n2645), .X($abc$9276$new_n2646)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11578 (
        .A($abc$9276$new_n1505), .B($abc$9276$new_n2640), .Y($abc$9276$new_n2647)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11579 (
        .A($abc$9276$new_n351), .B($abc$9276$new_n1504), .Y($abc$9276$new_n2648)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11580 (
        .A($abc$9276$new_n2647), .B($abc$9276$new_n2648), .Y($abc$9276$new_n2649)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11581 (
        .A($abc$9276$new_n2645), .B($abc$9276$new_n2649), .Y($abc$9276$new_n2650)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11582 (
        .A($abc$9276$new_n2646), .B($abc$9276$new_n2650), .Y($abc$9276$new_n2651)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11583 (
        .A($abc$9276$new_n378), .B($abc$9276$new_n2651), .X($abc$9276$new_n2652)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11584 (
        .A($abc$9276$new_n2652), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8979)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11585 (
        .A(CPU.I), .B($abc$9276$new_n742), .Y($abc$9276$new_n2654)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11586 (
        .A($abc$9276$new_n374), .B($abc$9276$new_n742), .X($abc$9276$new_n2655)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11587 (
        .A($abc$9276$new_n2654), .B($abc$9276$new_n2655), .Y($abc$9276$new_n2656)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11588 (
        .A($abc$9276$new_n1475), .B($abc$9276$new_n2656), .Y($abc$9276$new_n2657)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11589 (
        .A(oeb_16), .B(CPU.sei), .Y($abc$9276$new_n2658)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11590 (
        .A($abc$9276$new_n356), .B(CPU.I), .Y($abc$9276$new_n2659)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11591 (
        .A($abc$9276$new_n2658), .B($abc$9276$new_n2659), .Y($abc$9276$new_n2660)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11592 (
        .A($abc$9276$new_n355), .B($abc$9276$new_n2660), .Y($abc$9276$new_n2661)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11593 (
        .A(CPU.cli), .B(oeb_0), .Y($abc$9276$new_n2662)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11594 (
        .A($abc$9276$new_n2661), .B($abc$9276$new_n2662), .Y($abc$9276$new_n2663)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11595 (
        .A($abc$9276$new_n1476), .B($abc$9276$new_n2663), .Y($abc$9276$new_n2664)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11596 (
        .A($abc$9276$new_n2657), .B($abc$9276$new_n2664), .Y($abc$9276$new_n2665)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11597 (
        .A($abc$9276$new_n729), .B($abc$9276$new_n2665), .Y($abc$9276$new_n2666)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11598 (
        .A($abc$9276$new_n525), .B($abc$9276$new_n729), .X($abc$9276$new_n2667)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11599 (
        .A($abc$9276$new_n410), .B($abc$9276$new_n2667), .Y($abc$9276$new_n2668)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11600 (
        .A($abc$9276$new_n2668), .Y($abc$9276$new_n2669)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11601 (
        .A($abc$9276$new_n2666), .B($abc$9276$new_n2669), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8987)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11602 (
        .A($abc$9276$new_n1865), .B($abc$9276$new_n1916), .X($abc$9276$new_n2671)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11603 (
        .A(CPU.store), .B($abc$9276$new_n2671), .Y($abc$9276$new_n2672)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11604 (
        .A($abc$9276$new_n1352), .B($abc$9276$new_n2254), .X($abc$9276$new_n2673)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11605 (
        .A($abc$9276$new_n2673), .Y($abc$9276$new_n2674)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11606 (
        .A($abc$9276$new_n377), .B($abc$9276$new_n2671), .X($abc$9276$new_n2675)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11607 (
        .A($abc$9276$new_n2672), .B($abc$9276$new_n2675), .Y($abc$9276$new_n2676)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11608 (
        .A($abc$9276$new_n2673), .B($abc$9276$new_n2676), .X(out_32)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11609 (
        .A($abc$9276$new_n1436), .B($abc$9276$new_n2674), .Y($abc$9276$new_n2678)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11610 (
        .A($abc$9276$new_n353), .B($abc$9276$new_n385), .X($abc$9276$new_n2679)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11611 (
        .A($abc$9276$new_n1012), .B($abc$9276$new_n2679), .Y($abc$9276$new_n2680)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11612 (
        .A(CPU.C), .B($abc$9276$new_n2680), .Y($abc$9276$new_n2681)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11613 (
        .A(CPU.php), .B($abc$9276$new_n385), .X($abc$9276$new_n2682)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11614 (
        .A($abc$9276$new_n1351), .B($abc$9276$new_n2682), .Y($abc$9276$new_n2683)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11615 (
        .A(CPU.ADD), .B($abc$9276$new_n2683), .Y($abc$9276$new_n2684)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11616 (
        .A($abc$9276$new_n390), .B($abc$9276$new_n397), .Y($abc$9276$new_n2685)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11617 (
        .A(CPU.PC), .B($abc$9276$new_n2685), .Y($abc$9276$new_n2686)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11618 (
        .A(CPU.PC), .B($abc$9276$new_n1886), .Y($abc$9276$new_n2687)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11619 (
        .A($abc$9276$new_n2681), .B($abc$9276$new_n2687), .Y($abc$9276$new_n2688)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11620 (
        .A($abc$9276$new_n2684), .B($abc$9276$new_n2686), .Y($abc$9276$new_n2689)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11621 (
        .A($abc$9276$new_n2689), .Y($abc$9276$new_n2690)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11622 (
        .A($abc$9276$new_n2678), .B($abc$9276$new_n2690), .Y($abc$9276$new_n2691)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11623 (
        .A($abc$9276$new_n2688), .B($abc$9276$new_n2691), .X(out_24)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11624 (
        .A($abc$9276$new_n1521), .B($abc$9276$new_n2673), .X($abc$9276$new_n2693)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11625 (
        .A(CPU.ADD), .B($abc$9276$new_n2683), .Y($abc$9276$new_n2694)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11626 (
        .A($abc$9276$new_n2694), .Y($abc$9276$new_n2695)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11627 (
        .A(CPU.Z), .B($abc$9276$new_n2680), .Y($abc$9276$new_n2696)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11628 (
        .A(CPU.PC), .B($abc$9276$new_n2685), .Y($abc$9276$new_n2697)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11629 (
        .A(CPU.PC), .B($abc$9276$new_n1886), .Y($abc$9276$new_n2698)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11630 (
        .A($abc$9276$new_n2697), .B($abc$9276$new_n2698), .Y($abc$9276$new_n2699)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11631 (
        .A($abc$9276$new_n2699), .Y($abc$9276$new_n2700)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11632 (
        .A($abc$9276$new_n2696), .B($abc$9276$new_n2700), .Y($abc$9276$new_n2701)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11633 (
        .A($abc$9276$new_n2695), .B($abc$9276$new_n2701), .X($abc$9276$new_n2702)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11634 (
        .A($abc$9276$new_n2702), .Y($abc$9276$new_n2703)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11635 (
        .A($abc$9276$new_n2693), .B($abc$9276$new_n2703), .Y(out_25)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11636 (
        .A($abc$9276$new_n1544), .B($abc$9276$new_n2673), .X($abc$9276$new_n2705)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11637 (
        .A(CPU.I), .B($abc$9276$new_n2680), .Y($abc$9276$new_n2706)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11638 (
        .A($abc$9276$new_n2706), .Y($abc$9276$new_n2707)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11639 (
        .A(CPU.ADD), .B($abc$9276$new_n2683), .Y($abc$9276$new_n2708)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11640 (
        .A(CPU.PC), .B($abc$9276$new_n1886), .Y($abc$9276$new_n2709)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11641 (
        .A(CPU.PC), .B($abc$9276$new_n2685), .Y($abc$9276$new_n2710)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11642 (
        .A($abc$9276$new_n2709), .B($abc$9276$new_n2710), .Y($abc$9276$new_n2711)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11643 (
        .A($abc$9276$new_n2711), .Y($abc$9276$new_n2712)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11644 (
        .A($abc$9276$new_n2708), .B($abc$9276$new_n2712), .Y($abc$9276$new_n2713)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11645 (
        .A($abc$9276$new_n2707), .B($abc$9276$new_n2713), .X($abc$9276$new_n2714)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11646 (
        .A($abc$9276$new_n2714), .Y($abc$9276$new_n2715)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11647 (
        .A($abc$9276$new_n2705), .B($abc$9276$new_n2715), .Y(out_26)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11648 (
        .A($abc$9276$new_n1569), .B($abc$9276$new_n2673), .X($abc$9276$new_n2717)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11649 (
        .A(CPU.ADD), .B($abc$9276$new_n2683), .Y($abc$9276$new_n2718)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11650 (
        .A(CPU.D), .B($abc$9276$new_n2680), .Y($abc$9276$new_n2719)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11651 (
        .A(CPU.PC), .B($abc$9276$new_n2685), .Y($abc$9276$new_n2720)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11652 (
        .A(CPU.PC), .B($abc$9276$new_n1886), .Y($abc$9276$new_n2721)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11653 (
        .A($abc$9276$new_n2719), .B($abc$9276$new_n2721), .Y($abc$9276$new_n2722)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11654 (
        .A($abc$9276$new_n2718), .B($abc$9276$new_n2720), .Y($abc$9276$new_n2723)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11655 (
        .A($abc$9276$new_n2723), .Y($abc$9276$new_n2724)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11656 (
        .A($abc$9276$new_n2717), .B($abc$9276$new_n2724), .Y($abc$9276$new_n2725)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11657 (
        .A($abc$9276$new_n2722), .B($abc$9276$new_n2725), .X(out_27)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11658 (
        .A($abc$9276$new_n1595), .B($abc$9276$new_n2673), .X($abc$9276$new_n2727)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11659 (
        .A(CPU.ADD), .B($abc$9276$new_n2683), .Y($abc$9276$new_n2728)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11660 (
        .A($abc$9276$new_n2728), .Y($abc$9276$new_n2729)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11661 (
        .A(CPU.PC), .B($abc$9276$new_n2685), .Y($abc$9276$new_n2730)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11662 (
        .A(CPU.PC), .B($abc$9276$new_n1886), .Y($abc$9276$new_n2731)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11663 (
        .A($abc$9276$new_n2730), .B($abc$9276$new_n2731), .Y($abc$9276$new_n2732)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11664 (
        .A($abc$9276$new_n351), .B($abc$9276$new_n2679), .X($abc$9276$new_n2733)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11665 (
        .A($abc$9276$new_n757), .B($abc$9276$new_n1012), .X($abc$9276$new_n2734)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11666 (
        .A($abc$9276$new_n2733), .B($abc$9276$new_n2734), .Y($abc$9276$new_n2735)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11667 (
        .A($abc$9276$new_n2732), .B($abc$9276$new_n2735), .X($abc$9276$new_n2736)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11668 (
        .A($abc$9276$new_n2729), .B($abc$9276$new_n2736), .X($abc$9276$new_n2737)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11669 (
        .A($abc$9276$new_n2737), .Y($abc$9276$new_n2738)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11670 (
        .A($abc$9276$new_n2727), .B($abc$9276$new_n2738), .Y(out_28)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11671 (
        .A($abc$9276$new_n1621), .B($abc$9276$new_n2673), .X($abc$9276$new_n2740)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11672 (
        .A(CPU.ADD), .B($abc$9276$new_n2683), .Y($abc$9276$new_n2741)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11673 (
        .A($abc$9276$new_n2741), .Y($abc$9276$new_n2742)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11674 (
        .A($abc$9276$new_n1012), .B($abc$9276$new_n2733), .Y($abc$9276$new_n2743)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11675 (
        .A(CPU.PC), .B($abc$9276$new_n1886), .Y($abc$9276$new_n2744)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11676 (
        .A(CPU.PC), .B($abc$9276$new_n2685), .Y($abc$9276$new_n2745)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11677 (
        .A($abc$9276$new_n2744), .B($abc$9276$new_n2745), .Y($abc$9276$new_n2746)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11678 (
        .A($abc$9276$new_n2743), .B($abc$9276$new_n2746), .X($abc$9276$new_n2747)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11679 (
        .A($abc$9276$new_n2742), .B($abc$9276$new_n2747), .X($abc$9276$new_n2748)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11680 (
        .A($abc$9276$new_n2748), .Y($abc$9276$new_n2749)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11681 (
        .A($abc$9276$new_n2740), .B($abc$9276$new_n2749), .Y(out_29)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11682 (
        .A($abc$9276$new_n1647), .B($abc$9276$new_n2673), .X($abc$9276$new_n2751)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11683 (
        .A(CPU.ADD), .B($abc$9276$new_n2683), .Y($abc$9276$new_n2752)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11684 (
        .A(CPU.V), .B($abc$9276$new_n2680), .Y($abc$9276$new_n2753)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11685 (
        .A($abc$9276$new_n2753), .Y($abc$9276$new_n2754)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11686 (
        .A(CPU.PC), .B($abc$9276$new_n1886), .Y($abc$9276$new_n2755)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11687 (
        .A($abc$9276$new_n2755), .Y($abc$9276$new_n2756)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11688 (
        .A(CPU.PC), .B($abc$9276$new_n2685), .Y($abc$9276$new_n2757)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11689 (
        .A($abc$9276$new_n2752), .B($abc$9276$new_n2757), .Y($abc$9276$new_n2758)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11690 (
        .A($abc$9276$new_n2756), .B($abc$9276$new_n2758), .X($abc$9276$new_n2759)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11691 (
        .A($abc$9276$new_n2754), .B($abc$9276$new_n2759), .X($abc$9276$new_n2760)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11692 (
        .A($abc$9276$new_n2760), .Y($abc$9276$new_n2761)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11693 (
        .A($abc$9276$new_n2751), .B($abc$9276$new_n2761), .Y(out_30)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11694 (
        .A($abc$9276$new_n1673), .B($abc$9276$new_n2673), .X($abc$9276$new_n2763)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11695 (
        .A(CPU.N), .B($abc$9276$new_n2680), .Y($abc$9276$new_n2764)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11696 (
        .A($abc$9276$new_n2764), .Y($abc$9276$new_n2765)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11697 (
        .A($abc$9276$new_n372), .B($abc$9276$new_n2682), .X($abc$9276$new_n2766)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11698 (
        .A($abc$9276$new_n1358), .B($abc$9276$new_n2766), .Y($abc$9276$new_n2767)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11699 (
        .A(CPU.PC), .B($abc$9276$new_n2685), .Y($abc$9276$new_n2768)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11700 (
        .A(CPU.PC), .B($abc$9276$new_n1886), .Y($abc$9276$new_n2769)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11701 (
        .A($abc$9276$new_n2768), .B($abc$9276$new_n2769), .Y($abc$9276$new_n2770)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11702 (
        .A($abc$9276$new_n2767), .B($abc$9276$new_n2770), .X($abc$9276$new_n2771)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11703 (
        .A($abc$9276$new_n2765), .B($abc$9276$new_n2771), .X($abc$9276$new_n2772)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11704 (
        .A($abc$9276$new_n2772), .Y($abc$9276$new_n2773)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11705 (
        .A($abc$9276$new_n2763), .B($abc$9276$new_n2773), .Y(out_31)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11706 (
        .A(CPU.adc_sbc), .B(CPU.D), .Y($abc$9276$new_n2775)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$11707 (
        .A($abc$9276$new_n2775), .Y($abc$9276$flatten\CPU.$0\adj_bcd[0:0])
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9277 (
        .A(CPU.AXYS[3]), .Y($abc$9276$new_n346)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9278 (
        .A(CPU.AXYS[2]), .Y($abc$9276$new_n347)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9279 (
        .A(CPU.AXYS[0]), .Y($abc$9276$new_n348)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9280 (
        .A(CPU.V), .Y($abc$9276$new_n349)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9281 (
        .A(CPU.NMI_edge), .Y($abc$9276$new_n350)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9282 (
        .A(oeb_16), .Y($abc$9276$new_n351)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9283 (
        .A(CPU.plp), .Y($abc$9276$new_n352)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9284 (
        .A(CPU.php), .Y($abc$9276$new_n353)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9285 (
        .A(CPU.cld), .Y($abc$9276$new_n354)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9286 (
        .A(CPU.cli), .Y($abc$9276$new_n355)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9287 (
        .A(CPU.sei), .Y($abc$9276$new_n356)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9288 (
        .A(CPU.clv), .Y($abc$9276$new_n357)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9289 (
        .A(CPU.compare), .Y($abc$9276$new_n358)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9290 (
        .A(in_35), .Y($abc$9276$new_n359)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9291 (
        .A(CPU.cond_code), .Y($abc$9276$new_n360)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9292 (
        .A(CPU.N), .Y($abc$9276$new_n361)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9293 (
        .A(CPU.Z), .Y($abc$9276$new_n362)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9294 (
        .A(CPU.C), .Y($abc$9276$new_n363)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9295 (
        .A(CPU.IRHOLD), .Y($abc$9276$new_n364)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9296 (
        .A(CPU.IRHOLD), .Y($abc$9276$new_n365)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9297 (
        .A(CPU.IRHOLD), .Y($abc$9276$new_n366)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9298 (
        .A(CPU.IRHOLD), .Y($abc$9276$new_n367)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9299 (
        .A(CPU.IRHOLD), .Y($abc$9276$new_n368)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9300 (
        .A(CPU.IRHOLD), .Y($abc$9276$new_n369)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9301 (
        .A(CPU.IRHOLD), .Y($abc$9276$new_n370)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9302 (
        .A(CPU.src_reg), .Y($abc$9276$new_n371)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9303 (
        .A(CPU.ALU.N), .Y($abc$9276$new_n372)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9304 (
        .A(CPU.ADD), .Y($abc$9276$new_n373)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9305 (
        .A(CPU.ADD), .Y($abc$9276$new_n374)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9306 (
        .A(CPU.ADD), .Y($abc$9276$new_n375)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9307 (
        .A(CPU.ADD), .Y($abc$9276$new_n376)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9308 (
        .A(oeb_0), .Y($abc$9276$new_n377)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9309 (
        .A(rst_n), .Y($abc$9276$new_n378)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9310 (
        .A($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9180), .Y($abc$9276$new_n379)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9311 (
        .A(CPU.state), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9132), .X($abc$9276$new_n380)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9312 (
        .A($abc$9276$new_n380), .Y($abc$9276$new_n381)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9313 (
        .A(CPU.state), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9140), .X($abc$9276$new_n382)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9314 (
        .A(CPU.state), .B(CPU.state), .X($abc$9276$new_n383)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9315 (
        .A($abc$9276$new_n382), .B($abc$9276$new_n383), .X($abc$9276$new_n384)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9316 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n384), .X($abc$9276$new_n385)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9317 (
        .A(CPU.state), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9136), .X($abc$9276$new_n386)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9318 (
        .A($abc$9276$new_n382), .B($abc$9276$new_n386), .X($abc$9276$new_n387)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9319 (
        .A(CPU.state), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9134), .X($abc$9276$new_n388)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9320 (
        .A($abc$9276$new_n388), .Y($abc$9276$new_n389)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9321 (
        .A($abc$9276$new_n387), .B($abc$9276$new_n388), .X($abc$9276$new_n390)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9322 (
        .A($abc$9276$new_n390), .Y($abc$9276$new_n391)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9323 (
        .A($abc$9276$new_n385), .B($abc$9276$new_n390), .Y($abc$9276$new_n392)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9324 (
        .A(CPU.state), .B(CPU.state), .X($abc$9276$new_n393)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9325 (
        .A($abc$9276$new_n393), .Y($abc$9276$new_n394)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9326 (
        .A(CPU.state), .B(CPU.state), .X($abc$9276$new_n395)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9327 (
        .A($abc$9276$new_n386), .B($abc$9276$new_n395), .X($abc$9276$new_n396)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9328 (
        .A($abc$9276$new_n393), .B($abc$9276$new_n396), .X($abc$9276$new_n397)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9329 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n387), .X($abc$9276$new_n398)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9330 (
        .A(CPU.state), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9142), .X($abc$9276$new_n399)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9331 (
        .A(CPU.state), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9138), .X($abc$9276$new_n400)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9332 (
        .A($abc$9276$new_n399), .B($abc$9276$new_n400), .X($abc$9276$new_n401)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9333 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n401), .X($abc$9276$new_n402)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9334 (
        .A($abc$9276$new_n398), .B($abc$9276$new_n402), .Y($abc$9276$new_n403)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9335 (
        .A($abc$9276$new_n385), .B($abc$9276$new_n397), .Y($abc$9276$new_n404)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9336 (
        .A($abc$9276$new_n391), .B($abc$9276$new_n403), .X($abc$9276$new_n405)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9337 (
        .A($abc$9276$new_n404), .B($abc$9276$new_n405), .X($abc$9276$new_n406)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9338 (
        .A($abc$9276$new_n406), .Y($abc$9276$new_n407)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9339 (
        .A($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9142), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9140), .X($abc$9276$new_n408)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9340 (
        .A($abc$9276$new_n386), .B($abc$9276$new_n408), .X($abc$9276$new_n409)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9341 (
        .A($abc$9276$new_n393), .B($abc$9276$new_n409), .X($abc$9276$new_n410)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9342 (
        .A($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9138), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9136), .X($abc$9276$new_n411)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9343 (
        .A($abc$9276$new_n395), .B($abc$9276$new_n411), .X($abc$9276$new_n412)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9344 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n412), .X($abc$9276$new_n413)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9345 (
        .A($abc$9276$new_n410), .B($abc$9276$new_n413), .Y($abc$9276$new_n414)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9346 (
        .A($abc$9276$new_n408), .B($abc$9276$new_n411), .X($abc$9276$new_n415)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9347 (
        .A($abc$9276$new_n388), .B($abc$9276$new_n415), .X($abc$9276$new_n416)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9348 (
        .A($abc$9276$new_n416), .Y($abc$9276$new_n417)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9349 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n396), .X($abc$9276$new_n418)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9350 (
        .A($abc$9276$new_n416), .B($abc$9276$new_n418), .Y($abc$9276$new_n419)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9351 (
        .A($abc$9276$new_n382), .B($abc$9276$new_n411), .X($abc$9276$new_n420)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9352 (
        .A($abc$9276$new_n388), .B($abc$9276$new_n420), .X($abc$9276$new_n421)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9353 (
        .A($abc$9276$new_n421), .Y($abc$9276$new_n422)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9354 (
        .A($abc$9276$new_n388), .B($abc$9276$new_n412), .X($abc$9276$new_n423)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9355 (
        .A($abc$9276$new_n421), .B($abc$9276$new_n423), .Y($abc$9276$new_n424)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9356 (
        .A($abc$9276$new_n414), .B($abc$9276$new_n424), .X($abc$9276$new_n425)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9357 (
        .A($abc$9276$new_n419), .B($abc$9276$new_n425), .X($abc$9276$new_n426)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9358 (
        .A($abc$9276$new_n406), .B($abc$9276$new_n426), .X($abc$9276$new_n427)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9359 (
        .A($abc$9276$new_n393), .B($abc$9276$new_n412), .X($abc$9276$new_n428)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9360 (
        .A($abc$9276$new_n428), .Y($abc$9276$new_n429)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9361 (
        .A($abc$9276$new_n427), .B($abc$9276$new_n429), .X($abc$9276$new_n430)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9362 (
        .A($abc$9276$new_n383), .B($abc$9276$new_n395), .X($abc$9276$new_n431)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9363 (
        .A($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9134), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9132), .X($abc$9276$new_n432)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9364 (
        .A($abc$9276$new_n431), .B($abc$9276$new_n432), .X($abc$9276$new_n433)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9365 (
        .A($abc$9276$new_n383), .B($abc$9276$new_n408), .X($abc$9276$new_n434)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9366 (
        .A($abc$9276$new_n388), .B($abc$9276$new_n434), .X($abc$9276$new_n435)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9367 (
        .A($abc$9276$new_n433), .B($abc$9276$new_n435), .Y($abc$9276$new_n436)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9368 (
        .A($abc$9276$new_n393), .B($abc$9276$new_n420), .X($abc$9276$new_n437)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9369 (
        .A($abc$9276$new_n384), .B($abc$9276$new_n393), .X($abc$9276$new_n438)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9370 (
        .A($abc$9276$new_n437), .B($abc$9276$new_n438), .Y($abc$9276$new_n439)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9371 (
        .A($abc$9276$new_n436), .B($abc$9276$new_n439), .X($abc$9276$new_n440)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9372 (
        .A($abc$9276$new_n440), .Y($abc$9276$new_n441)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9373 (
        .A(CPU.src_reg), .B($abc$9276$new_n441), .Y($abc$9276$new_n442)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9374 (
        .A($abc$9276$new_n430), .B($abc$9276$new_n442), .X($abc$9276$new_n443)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9375 (
        .A(CPU.index_y), .B($abc$9276$new_n440), .Y($abc$9276$new_n444)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9376 (
        .A(CPU.dst_reg), .B($abc$9276$new_n429), .Y($abc$9276$new_n445)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9377 (
        .A($abc$9276$new_n444), .B($abc$9276$new_n445), .Y($abc$9276$new_n446)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9378 (
        .A($abc$9276$new_n427), .B($abc$9276$new_n446), .X($abc$9276$new_n447)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9379 (
        .A($abc$9276$new_n447), .Y($abc$9276$new_n448)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9380 (
        .A($abc$9276$new_n443), .B($abc$9276$new_n448), .Y($abc$9276$new_n449)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9381 (
        .A($abc$9276$new_n449), .Y($abc$9276$new_n450)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9382 (
        .A($abc$9276$new_n390), .B($abc$9276$new_n423), .Y($abc$9276$new_n451)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9383 (
        .A($abc$9276$new_n451), .Y($abc$9276$new_n452)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9384 (
        .A($abc$9276$new_n419), .B($abc$9276$new_n451), .X($abc$9276$new_n453)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9385 (
        .A(CPU.load_reg), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9226), .Y($abc$9276$new_n454)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9386 (
        .A($abc$9276$new_n428), .B($abc$9276$new_n454), .X($abc$9276$new_n455)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9387 (
        .A(oeb_0), .B($abc$9276$new_n428), .Y($abc$9276$new_n456)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9388 (
        .A($abc$9276$new_n455), .B($abc$9276$new_n456), .Y($abc$9276$new_n457)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9389 (
        .A($abc$9276$new_n453), .B($abc$9276$new_n457), .X($abc$9276$new_n458)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9390 (
        .A($abc$9276$new_n414), .B($abc$9276$new_n458), .X($abc$9276$new_n459)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9391 (
        .A(in_35), .B($abc$9276$new_n459), .Y($abc$9276$new_n460)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9392 (
        .A($abc$9276$new_n460), .Y($abc$9276$new_n461)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9393 (
        .A($abc$9276$new_n371), .B($abc$9276$new_n430), .X($abc$9276$new_n462)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9394 (
        .A(CPU.dst_reg), .B($abc$9276$new_n429), .Y($abc$9276$new_n463)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9395 (
        .A($abc$9276$new_n441), .B($abc$9276$new_n463), .Y($abc$9276$new_n464)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9396 (
        .A($abc$9276$new_n464), .Y($abc$9276$new_n465)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9397 (
        .A($abc$9276$new_n462), .B($abc$9276$new_n465), .Y($abc$9276$new_n466)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9398 (
        .A($abc$9276$new_n466), .Y($abc$9276$new_n467)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9399 (
        .A($abc$9276$new_n461), .B($abc$9276$new_n466), .Y($abc$9276$new_n468)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9400 (
        .A($abc$9276$new_n450), .B($abc$9276$new_n468), .X($abc$9276$new_n469)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9401 (
        .A($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9160), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9210), .X($abc$9276$new_n470)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9402 (
        .A($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9120), .B($abc$9276$new_n470), .X($abc$9276$new_n471)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9403 (
        .A(CPU.adc_bcd), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9160), .X($abc$9276$new_n472)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9404 (
        .A(CPU.ALU.HC), .B($abc$9276$new_n472), .X($abc$9276$new_n473)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9405 (
        .A($abc$9276$new_n471), .B($abc$9276$new_n473), .Y($abc$9276$new_n474)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9406 (
        .A(CPU.ALU.HC), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9210), .X($abc$9276$new_n475)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9407 (
        .A(CPU.adc_bcd), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9120), .X($abc$9276$new_n476)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9408 (
        .A($abc$9276$new_n475), .B($abc$9276$new_n476), .Y($abc$9276$new_n477)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9409 (
        .A($abc$9276$new_n474), .B($abc$9276$new_n477), .X($abc$9276$new_n478)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9410 (
        .A($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9160), .B($abc$9276$new_n478), .X($abc$9276$new_n479)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9411 (
        .A(oeb_0), .B($abc$9276$new_n479), .Y($abc$9276$new_n480)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9412 (
        .A($abc$9276$new_n373), .B($abc$9276$new_n480), .Y($abc$9276$new_n481)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9413 (
        .A($abc$9276$new_n373), .B($abc$9276$new_n480), .X($abc$9276$new_n482)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9414 (
        .A($abc$9276$new_n481), .B($abc$9276$new_n482), .Y($abc$9276$new_n483)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9415 (
        .A($abc$9276$new_n390), .B($abc$9276$new_n483), .Y($abc$9276$new_n484)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9416 (
        .A(in_35), .B(CPU.DIHOLD), .X($abc$9276$new_n485)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9417 (
        .A($abc$9276$new_n359), .B(in_16), .X($abc$9276$new_n486)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9418 (
        .A($abc$9276$new_n485), .B($abc$9276$new_n486), .Y($abc$9276$new_n487)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9419 (
        .A($abc$9276$new_n487), .Y(CPU.DIMUX)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9420 (
        .A($abc$9276$new_n390), .B(CPU.DIMUX), .X($abc$9276$new_n489)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9421 (
        .A($abc$9276$new_n489), .Y($abc$9276$new_n490)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9422 (
        .A($abc$9276$new_n461), .B($abc$9276$new_n484), .Y($abc$9276$new_n491)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9423 (
        .A($abc$9276$new_n490), .B($abc$9276$new_n491), .X($abc$9276$new_n492)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9424 (
        .A($abc$9276$new_n469), .B($abc$9276$new_n492), .X($abc$9276$new_n493)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9425 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n469), .Y($abc$9276$new_n494)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9426 (
        .A($abc$9276$new_n493), .B($abc$9276$new_n494), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8819)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9427 (
        .A(CPU.ADD), .B($abc$9276$new_n474), .Y($abc$9276$new_n496)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9428 (
        .A(CPU.ADD), .B($abc$9276$new_n474), .X($abc$9276$new_n497)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9429 (
        .A($abc$9276$new_n496), .B($abc$9276$new_n497), .Y($abc$9276$new_n498)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9430 (
        .A($abc$9276$new_n482), .B($abc$9276$new_n498), .Y($abc$9276$new_n499)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9431 (
        .A($abc$9276$new_n482), .B($abc$9276$new_n498), .X($abc$9276$new_n500)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9432 (
        .A($abc$9276$new_n499), .B($abc$9276$new_n500), .Y($abc$9276$new_n501)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9433 (
        .A($abc$9276$new_n390), .B($abc$9276$new_n501), .Y($abc$9276$new_n502)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9434 (
        .A(in_35), .B(CPU.DIHOLD), .X($abc$9276$new_n503)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9435 (
        .A($abc$9276$new_n359), .B(in_17), .X($abc$9276$new_n504)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9436 (
        .A($abc$9276$new_n503), .B($abc$9276$new_n504), .Y($abc$9276$new_n505)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9437 (
        .A($abc$9276$new_n505), .Y(CPU.DIMUX)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9438 (
        .A($abc$9276$new_n390), .B(CPU.DIMUX), .X($abc$9276$new_n507)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9439 (
        .A($abc$9276$new_n507), .Y($abc$9276$new_n508)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9440 (
        .A($abc$9276$new_n461), .B($abc$9276$new_n502), .Y($abc$9276$new_n509)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9441 (
        .A($abc$9276$new_n508), .B($abc$9276$new_n509), .X($abc$9276$new_n510)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9442 (
        .A($abc$9276$new_n469), .B($abc$9276$new_n510), .X($abc$9276$new_n511)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9443 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n469), .Y($abc$9276$new_n512)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9444 (
        .A($abc$9276$new_n511), .B($abc$9276$new_n512), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8821)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9445 (
        .A($abc$9276$new_n496), .B($abc$9276$new_n500), .Y($abc$9276$new_n514)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9446 (
        .A($abc$9276$new_n514), .Y($abc$9276$new_n515)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9447 (
        .A($abc$9276$new_n374), .B($abc$9276$new_n471), .X($abc$9276$new_n516)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9448 (
        .A($abc$9276$new_n374), .B($abc$9276$new_n471), .Y($abc$9276$new_n517)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9449 (
        .A($abc$9276$new_n516), .B($abc$9276$new_n517), .Y($abc$9276$new_n518)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9450 (
        .A($abc$9276$new_n515), .B($abc$9276$new_n518), .Y($abc$9276$new_n519)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9451 (
        .A($abc$9276$new_n515), .B($abc$9276$new_n518), .X($abc$9276$new_n520)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9452 (
        .A($abc$9276$new_n519), .B($abc$9276$new_n520), .Y($abc$9276$new_n521)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9453 (
        .A($abc$9276$new_n390), .B($abc$9276$new_n521), .Y($abc$9276$new_n522)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9454 (
        .A(in_35), .B(CPU.DIHOLD), .X($abc$9276$new_n523)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9455 (
        .A($abc$9276$new_n359), .B(in_18), .X($abc$9276$new_n524)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9456 (
        .A($abc$9276$new_n523), .B($abc$9276$new_n524), .Y($abc$9276$new_n525)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9457 (
        .A($abc$9276$new_n525), .Y(CPU.DIMUX)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9458 (
        .A($abc$9276$new_n390), .B(CPU.DIMUX), .X($abc$9276$new_n527)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9459 (
        .A($abc$9276$new_n461), .B($abc$9276$new_n527), .Y($abc$9276$new_n528)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9460 (
        .A($abc$9276$new_n528), .Y($abc$9276$new_n529)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9461 (
        .A($abc$9276$new_n522), .B($abc$9276$new_n529), .Y($abc$9276$new_n530)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9462 (
        .A($abc$9276$new_n469), .B($abc$9276$new_n530), .X($abc$9276$new_n531)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9463 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n469), .Y($abc$9276$new_n532)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9464 (
        .A($abc$9276$new_n531), .B($abc$9276$new_n532), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8823)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9465 (
        .A($abc$9276$new_n516), .B($abc$9276$new_n520), .Y($abc$9276$new_n534)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9466 (
        .A(CPU.ADD), .B($abc$9276$new_n473), .Y($abc$9276$new_n535)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9467 (
        .A(CPU.ADD), .B($abc$9276$new_n473), .X($abc$9276$new_n536)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9468 (
        .A($abc$9276$new_n535), .B($abc$9276$new_n536), .Y($abc$9276$new_n537)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9469 (
        .A($abc$9276$new_n537), .Y($abc$9276$new_n538)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9470 (
        .A($abc$9276$new_n534), .B($abc$9276$new_n538), .Y($abc$9276$new_n539)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9471 (
        .A($abc$9276$new_n534), .B($abc$9276$new_n538), .X($abc$9276$new_n540)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9472 (
        .A($abc$9276$new_n539), .B($abc$9276$new_n540), .Y($abc$9276$new_n541)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9473 (
        .A($abc$9276$new_n391), .B($abc$9276$new_n541), .X($abc$9276$new_n542)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9474 (
        .A(in_35), .B(CPU.DIHOLD), .X($abc$9276$new_n543)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9475 (
        .A($abc$9276$new_n359), .B(in_19), .X($abc$9276$new_n544)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9476 (
        .A($abc$9276$new_n543), .B($abc$9276$new_n544), .Y($abc$9276$new_n545)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9477 (
        .A($abc$9276$new_n545), .Y(CPU.DIMUX)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9478 (
        .A($abc$9276$new_n390), .B(CPU.DIMUX), .X($abc$9276$new_n547)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9479 (
        .A($abc$9276$new_n461), .B($abc$9276$new_n547), .Y($abc$9276$new_n548)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9480 (
        .A($abc$9276$new_n548), .Y($abc$9276$new_n549)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9481 (
        .A($abc$9276$new_n542), .B($abc$9276$new_n549), .Y($abc$9276$new_n550)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9482 (
        .A($abc$9276$new_n469), .B($abc$9276$new_n550), .X($abc$9276$new_n551)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9483 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n469), .Y($abc$9276$new_n552)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9484 (
        .A($abc$9276$new_n551), .B($abc$9276$new_n552), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8825)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9485 (
        .A($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9110), .B($abc$9276$new_n470), .X($abc$9276$new_n554)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9486 (
        .A(CPU.ALU.CO), .B($abc$9276$new_n472), .X($abc$9276$new_n555)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9487 (
        .A($abc$9276$new_n554), .B($abc$9276$new_n555), .Y($abc$9276$new_n556)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9488 (
        .A(CPU.ALU.CO), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9210), .X($abc$9276$new_n557)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9489 (
        .A(CPU.adc_bcd), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9110), .X($abc$9276$new_n558)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9490 (
        .A($abc$9276$new_n557), .B($abc$9276$new_n558), .Y($abc$9276$new_n559)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9491 (
        .A($abc$9276$new_n556), .B($abc$9276$new_n559), .X($abc$9276$new_n560)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9492 (
        .A($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9160), .B($abc$9276$new_n560), .X($abc$9276$new_n561)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9493 (
        .A(oeb_0), .B($abc$9276$new_n561), .Y($abc$9276$new_n562)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9494 (
        .A($abc$9276$new_n375), .B($abc$9276$new_n562), .Y($abc$9276$new_n563)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9495 (
        .A($abc$9276$new_n375), .B($abc$9276$new_n562), .X($abc$9276$new_n564)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9496 (
        .A($abc$9276$new_n563), .B($abc$9276$new_n564), .Y($abc$9276$new_n565)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9497 (
        .A($abc$9276$new_n390), .B($abc$9276$new_n565), .Y($abc$9276$new_n566)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9498 (
        .A(in_35), .B(in_20), .Y($abc$9276$new_n567)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9499 (
        .A($abc$9276$new_n359), .B(CPU.DIHOLD), .Y($abc$9276$new_n568)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9500 (
        .A($abc$9276$new_n567), .B($abc$9276$new_n568), .Y(CPU.DIMUX)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9501 (
        .A($abc$9276$new_n390), .B(CPU.DIMUX), .X($abc$9276$new_n570)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9502 (
        .A($abc$9276$new_n570), .Y($abc$9276$new_n571)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9503 (
        .A($abc$9276$new_n461), .B($abc$9276$new_n566), .Y($abc$9276$new_n572)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9504 (
        .A($abc$9276$new_n571), .B($abc$9276$new_n572), .X($abc$9276$new_n573)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9505 (
        .A($abc$9276$new_n469), .B($abc$9276$new_n573), .X($abc$9276$new_n574)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9506 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n469), .Y($abc$9276$new_n575)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9507 (
        .A($abc$9276$new_n574), .B($abc$9276$new_n575), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8827)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9508 (
        .A(CPU.ADD), .B($abc$9276$new_n556), .Y($abc$9276$new_n577)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9509 (
        .A(CPU.ADD), .B($abc$9276$new_n556), .X($abc$9276$new_n578)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9510 (
        .A($abc$9276$new_n577), .B($abc$9276$new_n578), .Y($abc$9276$new_n579)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9511 (
        .A($abc$9276$new_n564), .B($abc$9276$new_n579), .Y($abc$9276$new_n580)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9512 (
        .A($abc$9276$new_n564), .B($abc$9276$new_n579), .X($abc$9276$new_n581)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9513 (
        .A($abc$9276$new_n580), .B($abc$9276$new_n581), .Y($abc$9276$new_n582)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9514 (
        .A($abc$9276$new_n390), .B($abc$9276$new_n582), .Y($abc$9276$new_n583)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9515 (
        .A(in_35), .B(CPU.DIHOLD), .X($abc$9276$new_n584)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9516 (
        .A($abc$9276$new_n359), .B(in_21), .X($abc$9276$new_n585)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9517 (
        .A($abc$9276$new_n584), .B($abc$9276$new_n585), .Y($abc$9276$new_n586)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9518 (
        .A($abc$9276$new_n586), .Y(CPU.DIMUX)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9519 (
        .A($abc$9276$new_n390), .B(CPU.DIMUX), .X($abc$9276$new_n588)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9520 (
        .A($abc$9276$new_n588), .Y($abc$9276$new_n589)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9521 (
        .A($abc$9276$new_n461), .B($abc$9276$new_n583), .Y($abc$9276$new_n590)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9522 (
        .A($abc$9276$new_n589), .B($abc$9276$new_n590), .X($abc$9276$new_n591)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9523 (
        .A($abc$9276$new_n469), .B($abc$9276$new_n591), .X($abc$9276$new_n592)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9524 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n469), .Y($abc$9276$new_n593)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9525 (
        .A($abc$9276$new_n592), .B($abc$9276$new_n593), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8829)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9526 (
        .A($abc$9276$new_n577), .B($abc$9276$new_n581), .Y($abc$9276$new_n595)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9527 (
        .A($abc$9276$new_n595), .Y($abc$9276$new_n596)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9528 (
        .A($abc$9276$new_n376), .B($abc$9276$new_n554), .X($abc$9276$new_n597)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9529 (
        .A($abc$9276$new_n376), .B($abc$9276$new_n554), .Y($abc$9276$new_n598)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9530 (
        .A($abc$9276$new_n597), .B($abc$9276$new_n598), .Y($abc$9276$new_n599)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9531 (
        .A($abc$9276$new_n596), .B($abc$9276$new_n599), .Y($abc$9276$new_n600)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9532 (
        .A($abc$9276$new_n596), .B($abc$9276$new_n599), .X($abc$9276$new_n601)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9533 (
        .A($abc$9276$new_n600), .B($abc$9276$new_n601), .Y($abc$9276$new_n602)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9534 (
        .A($abc$9276$new_n390), .B($abc$9276$new_n602), .Y($abc$9276$new_n603)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9535 (
        .A(in_35), .B(CPU.DIHOLD), .X($abc$9276$new_n604)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9536 (
        .A($abc$9276$new_n359), .B(in_22), .X($abc$9276$new_n605)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9537 (
        .A($abc$9276$new_n604), .B($abc$9276$new_n605), .Y($abc$9276$new_n606)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9538 (
        .A($abc$9276$new_n606), .Y(CPU.DIMUX)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9539 (
        .A($abc$9276$new_n390), .B(CPU.DIMUX), .X($abc$9276$new_n608)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9540 (
        .A($abc$9276$new_n461), .B($abc$9276$new_n608), .Y($abc$9276$new_n609)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9541 (
        .A($abc$9276$new_n609), .Y($abc$9276$new_n610)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9542 (
        .A($abc$9276$new_n603), .B($abc$9276$new_n610), .Y($abc$9276$new_n611)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9543 (
        .A($abc$9276$new_n469), .B($abc$9276$new_n611), .X($abc$9276$new_n612)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9544 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n469), .Y($abc$9276$new_n613)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9545 (
        .A($abc$9276$new_n612), .B($abc$9276$new_n613), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8831)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9546 (
        .A($abc$9276$new_n597), .B($abc$9276$new_n601), .Y($abc$9276$new_n615)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9547 (
        .A(CPU.ALU.N), .B($abc$9276$new_n555), .Y($abc$9276$new_n616)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9548 (
        .A(CPU.ALU.N), .B($abc$9276$new_n555), .X($abc$9276$new_n617)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9549 (
        .A($abc$9276$new_n616), .B($abc$9276$new_n617), .Y($abc$9276$new_n618)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9550 (
        .A($abc$9276$new_n615), .B($abc$9276$new_n618), .X($abc$9276$new_n619)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9551 (
        .A($abc$9276$new_n615), .B($abc$9276$new_n618), .Y($abc$9276$new_n620)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9552 (
        .A($abc$9276$new_n619), .B($abc$9276$new_n620), .Y($abc$9276$new_n621)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9553 (
        .A($abc$9276$new_n390), .B($abc$9276$new_n621), .Y($abc$9276$new_n622)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9554 (
        .A($abc$9276$new_n359), .B(CPU.DIHOLD), .Y($abc$9276$new_n623)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9555 (
        .A(in_35), .B(in_23), .Y($abc$9276$new_n624)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9556 (
        .A($abc$9276$new_n623), .B($abc$9276$new_n624), .Y(CPU.DIMUX)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9557 (
        .A($abc$9276$new_n390), .B(CPU.DIMUX), .X($abc$9276$new_n626)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9558 (
        .A($abc$9276$new_n461), .B($abc$9276$new_n626), .Y($abc$9276$new_n627)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9559 (
        .A($abc$9276$new_n627), .Y($abc$9276$new_n628)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9560 (
        .A($abc$9276$new_n622), .B($abc$9276$new_n628), .Y($abc$9276$new_n629)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9561 (
        .A($abc$9276$new_n469), .B($abc$9276$new_n629), .X($abc$9276$new_n630)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9562 (
        .A(CPU.AXYS[3]), .B($abc$9276$new_n469), .Y($abc$9276$new_n631)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9563 (
        .A($abc$9276$new_n630), .B($abc$9276$new_n631), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8833)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9564 (
        .A($abc$9276$new_n449), .B($abc$9276$new_n468), .X($abc$9276$new_n633)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9565 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n633), .Y($abc$9276$new_n634)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9566 (
        .A($abc$9276$new_n492), .B($abc$9276$new_n633), .X($abc$9276$new_n635)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9567 (
        .A($abc$9276$new_n634), .B($abc$9276$new_n635), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8835)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9568 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n633), .Y($abc$9276$new_n637)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9569 (
        .A($abc$9276$new_n510), .B($abc$9276$new_n633), .X($abc$9276$new_n638)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9570 (
        .A($abc$9276$new_n637), .B($abc$9276$new_n638), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8837)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9571 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n633), .Y($abc$9276$new_n640)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9572 (
        .A($abc$9276$new_n530), .B($abc$9276$new_n633), .X($abc$9276$new_n641)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9573 (
        .A($abc$9276$new_n640), .B($abc$9276$new_n641), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8839)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9574 (
        .A($abc$9276$new_n550), .B($abc$9276$new_n633), .X($abc$9276$new_n643)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9575 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n633), .Y($abc$9276$new_n644)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9576 (
        .A($abc$9276$new_n643), .B($abc$9276$new_n644), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8841)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9577 (
        .A($abc$9276$new_n573), .B($abc$9276$new_n633), .X($abc$9276$new_n646)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9578 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n633), .Y($abc$9276$new_n647)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9579 (
        .A($abc$9276$new_n646), .B($abc$9276$new_n647), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8843)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9580 (
        .A($abc$9276$new_n591), .B($abc$9276$new_n633), .X($abc$9276$new_n649)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9581 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n633), .Y($abc$9276$new_n650)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9582 (
        .A($abc$9276$new_n649), .B($abc$9276$new_n650), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8845)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9583 (
        .A($abc$9276$new_n611), .B($abc$9276$new_n633), .X($abc$9276$new_n652)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9584 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n633), .Y($abc$9276$new_n653)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9585 (
        .A($abc$9276$new_n652), .B($abc$9276$new_n653), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8847)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9586 (
        .A(CPU.AXYS[2]), .B($abc$9276$new_n633), .Y($abc$9276$new_n655)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9587 (
        .A($abc$9276$new_n629), .B($abc$9276$new_n633), .X($abc$9276$new_n656)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9588 (
        .A($abc$9276$new_n655), .B($abc$9276$new_n656), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8849)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9589 (
        .A($abc$9276$new_n449), .B($abc$9276$new_n467), .Y($abc$9276$new_n658)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9590 (
        .A($abc$9276$new_n460), .B($abc$9276$new_n658), .X($abc$9276$new_n659)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9591 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n659), .Y($abc$9276$new_n660)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9592 (
        .A($abc$9276$new_n492), .B($abc$9276$new_n659), .X($abc$9276$new_n661)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9593 (
        .A($abc$9276$new_n660), .B($abc$9276$new_n661), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8851)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9594 (
        .A($abc$9276$new_n510), .B($abc$9276$new_n659), .X($abc$9276$new_n663)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9595 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n659), .Y($abc$9276$new_n664)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9596 (
        .A($abc$9276$new_n663), .B($abc$9276$new_n664), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8853)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9597 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n659), .Y($abc$9276$new_n666)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9598 (
        .A($abc$9276$new_n530), .B($abc$9276$new_n659), .X($abc$9276$new_n667)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9599 (
        .A($abc$9276$new_n666), .B($abc$9276$new_n667), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8855)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9600 (
        .A($abc$9276$new_n550), .B($abc$9276$new_n659), .X($abc$9276$new_n669)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9601 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n659), .Y($abc$9276$new_n670)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9602 (
        .A($abc$9276$new_n669), .B($abc$9276$new_n670), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8857)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9603 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n659), .Y($abc$9276$new_n672)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9604 (
        .A($abc$9276$new_n573), .B($abc$9276$new_n659), .X($abc$9276$new_n673)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9605 (
        .A($abc$9276$new_n672), .B($abc$9276$new_n673), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8859)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9606 (
        .A($abc$9276$new_n591), .B($abc$9276$new_n659), .X($abc$9276$new_n675)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9607 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n659), .Y($abc$9276$new_n676)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9608 (
        .A($abc$9276$new_n675), .B($abc$9276$new_n676), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8861)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9609 (
        .A($abc$9276$new_n611), .B($abc$9276$new_n659), .X($abc$9276$new_n678)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9610 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n659), .Y($abc$9276$new_n679)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9611 (
        .A($abc$9276$new_n678), .B($abc$9276$new_n679), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8863)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9612 (
        .A($abc$9276$new_n629), .B($abc$9276$new_n659), .X($abc$9276$new_n681)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9613 (
        .A(CPU.AXYS[1]), .B($abc$9276$new_n659), .Y($abc$9276$new_n682)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9614 (
        .A($abc$9276$new_n681), .B($abc$9276$new_n682), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8865)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9615 (
        .A($abc$9276$new_n449), .B($abc$9276$new_n466), .X($abc$9276$new_n684)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9616 (
        .A($abc$9276$new_n460), .B($abc$9276$new_n684), .X($abc$9276$new_n685)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9617 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n685), .Y($abc$9276$new_n686)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9618 (
        .A($abc$9276$new_n492), .B($abc$9276$new_n685), .X($abc$9276$new_n687)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9619 (
        .A($abc$9276$new_n686), .B($abc$9276$new_n687), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8867)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9620 (
        .A($abc$9276$new_n510), .B($abc$9276$new_n685), .X($abc$9276$new_n689)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9621 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n685), .Y($abc$9276$new_n690)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9622 (
        .A($abc$9276$new_n689), .B($abc$9276$new_n690), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8869)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9623 (
        .A($abc$9276$new_n530), .B($abc$9276$new_n685), .X($abc$9276$new_n692)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9624 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n685), .Y($abc$9276$new_n693)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9625 (
        .A($abc$9276$new_n692), .B($abc$9276$new_n693), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8871)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9626 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n685), .Y($abc$9276$new_n695)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9627 (
        .A($abc$9276$new_n550), .B($abc$9276$new_n685), .X($abc$9276$new_n696)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9628 (
        .A($abc$9276$new_n695), .B($abc$9276$new_n696), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8873)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9629 (
        .A($abc$9276$new_n573), .B($abc$9276$new_n685), .X($abc$9276$new_n698)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9630 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n685), .Y($abc$9276$new_n699)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9631 (
        .A($abc$9276$new_n698), .B($abc$9276$new_n699), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8875)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9632 (
        .A($abc$9276$new_n591), .B($abc$9276$new_n685), .X($abc$9276$new_n701)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9633 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n685), .Y($abc$9276$new_n702)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9634 (
        .A($abc$9276$new_n701), .B($abc$9276$new_n702), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8877)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9635 (
        .A($abc$9276$new_n611), .B($abc$9276$new_n685), .X($abc$9276$new_n704)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9636 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n685), .Y($abc$9276$new_n705)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9637 (
        .A($abc$9276$new_n704), .B($abc$9276$new_n705), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8879)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9638 (
        .A(CPU.AXYS[0]), .B($abc$9276$new_n685), .Y($abc$9276$new_n707)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9639 (
        .A($abc$9276$new_n629), .B($abc$9276$new_n685), .X($abc$9276$new_n708)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9640 (
        .A($abc$9276$new_n707), .B($abc$9276$new_n708), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8881)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9641 (
        .A(CPU.ALU.AI7), .B(CPU.ALU.CO), .X($abc$9276$new_n710)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9642 (
        .A(CPU.ALU.AI7), .B(CPU.ALU.CO), .Y($abc$9276$new_n711)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9643 (
        .A($abc$9276$new_n710), .B($abc$9276$new_n711), .Y($abc$9276$new_n712)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9644 (
        .A(CPU.ALU.BI7), .B(CPU.ALU.N), .Y($abc$9276$new_n713)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9645 (
        .A(CPU.ALU.BI7), .B(CPU.ALU.N), .X($abc$9276$new_n714)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9646 (
        .A($abc$9276$new_n713), .B($abc$9276$new_n714), .Y($abc$9276$new_n715)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9647 (
        .A($abc$9276$new_n712), .B($abc$9276$new_n715), .Y($abc$9276$new_n716)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9648 (
        .A($abc$9276$new_n712), .B($abc$9276$new_n715), .X($abc$9276$new_n717)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9649 (
        .A($abc$9276$new_n716), .B($abc$9276$new_n717), .Y($abc$9276$new_n718)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9650 (
        .A($abc$9276$new_n357), .B(CPU.adc_sbc), .Y($abc$9276$new_n719)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9651 (
        .A($abc$9276$new_n719), .Y($abc$9276$new_n720)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9652 (
        .A($abc$9276$new_n718), .B($abc$9276$new_n720), .Y($abc$9276$new_n721)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9653 (
        .A(CPU.clv), .B($abc$9276$new_n377), .Y($abc$9276$new_n722)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9654 (
        .A($abc$9276$new_n352), .B($abc$9276$new_n722), .Y($abc$9276$new_n723)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9655 (
        .A($abc$9276$new_n723), .Y($abc$9276$new_n724)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9656 (
        .A($abc$9276$new_n721), .B($abc$9276$new_n724), .Y($abc$9276$new_n725)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9657 (
        .A($abc$9276$new_n725), .Y($abc$9276$new_n726)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9658 (
        .A(CPU.plp), .B(CPU.ADD), .Y($abc$9276$new_n727)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9659 (
        .A($abc$9276$new_n400), .B($abc$9276$new_n408), .X($abc$9276$new_n728)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9660 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n728), .X($abc$9276$new_n729)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9661 (
        .A($abc$9276$new_n729), .Y($abc$9276$new_n730)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9662 (
        .A($abc$9276$new_n429), .B($abc$9276$new_n729), .Y($abc$9276$new_n731)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9663 (
        .A($abc$9276$new_n731), .Y($abc$9276$new_n732)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9664 (
        .A($abc$9276$new_n727), .B($abc$9276$new_n732), .Y($abc$9276$new_n733)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9665 (
        .A($abc$9276$new_n726), .B($abc$9276$new_n733), .X($abc$9276$new_n734)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9666 (
        .A($abc$9276$new_n399), .B($abc$9276$new_n411), .X($abc$9276$new_n735)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9667 (
        .A($abc$9276$new_n393), .B($abc$9276$new_n735), .X($abc$9276$new_n736)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9668 (
        .A($abc$9276$new_n736), .Y($abc$9276$new_n737)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9669 (
        .A(CPU.bit_ins), .B($abc$9276$new_n737), .Y($abc$9276$new_n738)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9670 (
        .A($abc$9276$new_n429), .B($abc$9276$new_n738), .X($abc$9276$new_n739)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9671 (
        .A($abc$9276$new_n729), .B($abc$9276$new_n739), .Y($abc$9276$new_n740)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9672 (
        .A($abc$9276$new_n740), .Y($abc$9276$new_n741)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9673 (
        .A($abc$9276$new_n352), .B($abc$9276$new_n428), .X($abc$9276$new_n742)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9674 (
        .A(CPU.clv), .B(CPU.adc_sbc), .X($abc$9276$new_n743)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9675 (
        .A(CPU.plp), .B($abc$9276$new_n743), .X($abc$9276$new_n744)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9676 (
        .A($abc$9276$new_n429), .B($abc$9276$new_n744), .Y($abc$9276$new_n745)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9677 (
        .A($abc$9276$new_n349), .B($abc$9276$new_n745), .Y($abc$9276$new_n746)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9678 (
        .A($abc$9276$new_n741), .B($abc$9276$new_n746), .Y($abc$9276$new_n747)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9679 (
        .A(CPU.DIMUX), .B($abc$9276$new_n740), .Y($abc$9276$new_n748)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9680 (
        .A($abc$9276$new_n747), .B($abc$9276$new_n748), .Y($abc$9276$new_n749)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9681 (
        .A($abc$9276$new_n734), .B($abc$9276$new_n749), .Y($abc$9276$new_n750)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9682 (
        .A($abc$9276$new_n750), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8883)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9683 (
        .A($abc$9276$new_n359), .B($abc$9276$new_n428), .X($abc$9276$new_n752)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9684 (
        .A($abc$9276$new_n752), .Y($abc$9276$new_n753)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9685 (
        .A(CPU.plp), .B($abc$9276$new_n752), .Y($abc$9276$new_n754)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9686 (
        .A(CPU.IRHOLD_valid), .B(CPU.DIMUX), .X($abc$9276$new_n755)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9687 (
        .A(in_33), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9174), .Y($abc$9276$new_n756)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9688 (
        .A(CPU.NMI_edge), .B(in_33), .X($abc$9276$new_n757)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9689 (
        .A(CPU.NMI_edge), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9174), .X($abc$9276$new_n758)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9690 (
        .A($abc$9276$new_n757), .B($abc$9276$new_n758), .Y($abc$9276$new_n759)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9691 (
        .A($abc$9276$new_n350), .B($abc$9276$new_n756), .Y($abc$9276$new_n760)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9692 (
        .A(CPU.IRHOLD_valid), .B($abc$9276$new_n369), .Y($abc$9276$new_n761)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9693 (
        .A($abc$9276$new_n755), .B($abc$9276$new_n761), .Y($abc$9276$new_n762)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9694 (
        .A($abc$9276$new_n760), .B($abc$9276$new_n762), .X($abc$9276$new_n763)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9695 (
        .A($abc$9276$new_n763), .Y($abc$9276$new_n764)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9696 (
        .A(CPU.IRHOLD_valid), .B(CPU.DIMUX), .X($abc$9276$new_n765)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9697 (
        .A(CPU.IRHOLD_valid), .B($abc$9276$new_n370), .Y($abc$9276$new_n766)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9698 (
        .A($abc$9276$new_n759), .B($abc$9276$new_n766), .Y($abc$9276$new_n767)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9699 (
        .A($abc$9276$new_n767), .Y($abc$9276$new_n768)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9700 (
        .A($abc$9276$new_n765), .B($abc$9276$new_n768), .Y($abc$9276$new_n769)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9701 (
        .A($abc$9276$new_n769), .Y($abc$9276$new_n770)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9702 (
        .A(CPU.IRHOLD_valid), .B(CPU.DIMUX), .X($abc$9276$new_n771)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9703 (
        .A(CPU.IRHOLD_valid), .B($abc$9276$new_n368), .Y($abc$9276$new_n772)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9704 (
        .A($abc$9276$new_n771), .B($abc$9276$new_n772), .Y($abc$9276$new_n773)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9705 (
        .A($abc$9276$new_n760), .B($abc$9276$new_n773), .X($abc$9276$new_n774)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9706 (
        .A($abc$9276$new_n774), .Y($abc$9276$new_n775)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9707 (
        .A(oeb_0), .B($abc$9276$new_n760), .Y($abc$9276$new_n776)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9708 (
        .A($abc$9276$new_n774), .B($abc$9276$new_n776), .Y($abc$9276$new_n777)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9709 (
        .A($abc$9276$new_n777), .Y($abc$9276$new_n778)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9710 (
        .A($abc$9276$new_n769), .B($abc$9276$new_n776), .Y($abc$9276$new_n779)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9711 (
        .A($abc$9276$new_n779), .Y($abc$9276$new_n780)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9712 (
        .A($abc$9276$new_n774), .B($abc$9276$new_n780), .Y($abc$9276$new_n781)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9713 (
        .A($abc$9276$new_n781), .Y($abc$9276$new_n782)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9714 (
        .A(CPU.IRHOLD_valid), .B($abc$9276$new_n586), .X($abc$9276$new_n783)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9715 (
        .A(CPU.IRHOLD_valid), .B(CPU.IRHOLD), .Y($abc$9276$new_n784)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9716 (
        .A($abc$9276$new_n783), .B($abc$9276$new_n784), .Y($abc$9276$new_n785)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9717 (
        .A($abc$9276$new_n759), .B($abc$9276$new_n785), .Y($abc$9276$new_n786)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9718 (
        .A($abc$9276$new_n777), .B($abc$9276$new_n786), .X($abc$9276$new_n787)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9719 (
        .A($abc$9276$new_n781), .B($abc$9276$new_n786), .X($abc$9276$new_n788)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9720 (
        .A($abc$9276$new_n763), .B($abc$9276$new_n776), .Y($abc$9276$new_n789)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9721 (
        .A($abc$9276$new_n788), .B($abc$9276$new_n789), .X($abc$9276$new_n790)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9722 (
        .A(CPU.IRHOLD_valid), .B(CPU.DIMUX), .X($abc$9276$new_n791)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9723 (
        .A(CPU.IRHOLD_valid), .B($abc$9276$new_n365), .Y($abc$9276$new_n792)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9724 (
        .A($abc$9276$new_n759), .B($abc$9276$new_n792), .Y($abc$9276$new_n793)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9725 (
        .A($abc$9276$new_n793), .Y($abc$9276$new_n794)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9726 (
        .A($abc$9276$new_n791), .B($abc$9276$new_n794), .Y($abc$9276$new_n795)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9727 (
        .A($abc$9276$new_n795), .Y($abc$9276$new_n796)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9728 (
        .A(CPU.IRHOLD_valid), .B(CPU.DIMUX), .X($abc$9276$new_n797)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9729 (
        .A(CPU.IRHOLD_valid), .B($abc$9276$new_n364), .Y($abc$9276$new_n798)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9730 (
        .A($abc$9276$new_n797), .B($abc$9276$new_n798), .Y($abc$9276$new_n799)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9731 (
        .A($abc$9276$new_n760), .B($abc$9276$new_n799), .X($abc$9276$new_n800)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9732 (
        .A($abc$9276$new_n800), .Y($abc$9276$new_n801)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9733 (
        .A($abc$9276$new_n776), .B($abc$9276$new_n800), .Y($abc$9276$new_n802)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9734 (
        .A($abc$9276$new_n796), .B($abc$9276$new_n802), .X($abc$9276$new_n803)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9735 (
        .A($abc$9276$new_n803), .Y($abc$9276$new_n804)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9736 (
        .A(CPU.IRHOLD_valid), .B(CPU.DIMUX), .X($abc$9276$new_n805)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9737 (
        .A(CPU.IRHOLD_valid), .B($abc$9276$new_n367), .Y($abc$9276$new_n806)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9738 (
        .A($abc$9276$new_n805), .B($abc$9276$new_n806), .Y($abc$9276$new_n807)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9739 (
        .A($abc$9276$new_n760), .B($abc$9276$new_n807), .X($abc$9276$new_n808)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9740 (
        .A(CPU.IRHOLD_valid), .B(CPU.DIMUX), .X($abc$9276$new_n809)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9741 (
        .A(CPU.IRHOLD_valid), .B($abc$9276$new_n366), .Y($abc$9276$new_n810)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9742 (
        .A($abc$9276$new_n759), .B($abc$9276$new_n810), .Y($abc$9276$new_n811)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9743 (
        .A($abc$9276$new_n811), .Y($abc$9276$new_n812)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9744 (
        .A($abc$9276$new_n809), .B($abc$9276$new_n812), .Y($abc$9276$new_n813)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9745 (
        .A($abc$9276$new_n776), .B($abc$9276$new_n813), .Y($abc$9276$new_n814)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9746 (
        .A($abc$9276$new_n808), .B($abc$9276$new_n814), .X($abc$9276$new_n815)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9747 (
        .A($abc$9276$new_n803), .B($abc$9276$new_n815), .X($abc$9276$new_n816)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9748 (
        .A($abc$9276$new_n752), .B($abc$9276$new_n816), .X($abc$9276$new_n817)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9749 (
        .A($abc$9276$new_n790), .B($abc$9276$new_n817), .X($abc$9276$new_n818)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9750 (
        .A($abc$9276$new_n754), .B($abc$9276$new_n818), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8889)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9751 (
        .A(CPU.php), .B($abc$9276$new_n752), .Y($abc$9276$new_n820)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9752 (
        .A($abc$9276$new_n782), .B($abc$9276$new_n786), .Y($abc$9276$new_n821)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9753 (
        .A($abc$9276$new_n764), .B($abc$9276$new_n821), .X($abc$9276$new_n822)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9754 (
        .A($abc$9276$new_n817), .B($abc$9276$new_n822), .X($abc$9276$new_n823)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9755 (
        .A($abc$9276$new_n820), .B($abc$9276$new_n823), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8891)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9756 (
        .A(CPU.clc), .B($abc$9276$new_n752), .Y($abc$9276$new_n825)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9757 (
        .A($abc$9276$new_n763), .B($abc$9276$new_n780), .Y($abc$9276$new_n826)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9758 (
        .A($abc$9276$new_n776), .B($abc$9276$new_n786), .Y($abc$9276$new_n827)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9759 (
        .A($abc$9276$new_n827), .Y($abc$9276$new_n828)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9760 (
        .A($abc$9276$new_n774), .B($abc$9276$new_n827), .X($abc$9276$new_n829)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9761 (
        .A($abc$9276$new_n817), .B($abc$9276$new_n829), .X($abc$9276$new_n830)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9762 (
        .A($abc$9276$new_n826), .B($abc$9276$new_n830), .X($abc$9276$new_n831)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9763 (
        .A($abc$9276$new_n825), .B($abc$9276$new_n831), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8893)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9764 (
        .A(CPU.sec), .B($abc$9276$new_n752), .Y($abc$9276$new_n833)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9765 (
        .A($abc$9276$new_n777), .B($abc$9276$new_n827), .Y($abc$9276$new_n834)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9766 (
        .A($abc$9276$new_n817), .B($abc$9276$new_n834), .X($abc$9276$new_n835)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9767 (
        .A($abc$9276$new_n826), .B($abc$9276$new_n835), .X($abc$9276$new_n836)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9768 (
        .A($abc$9276$new_n833), .B($abc$9276$new_n836), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8895)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9769 (
        .A(CPU.cld), .B($abc$9276$new_n752), .Y($abc$9276$new_n838)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9770 (
        .A($abc$9276$new_n779), .B($abc$9276$new_n789), .Y($abc$9276$new_n839)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9771 (
        .A($abc$9276$new_n830), .B($abc$9276$new_n839), .X($abc$9276$new_n840)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9772 (
        .A($abc$9276$new_n838), .B($abc$9276$new_n840), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8897)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9773 (
        .A(CPU.sed), .B($abc$9276$new_n752), .Y($abc$9276$new_n842)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9774 (
        .A($abc$9276$new_n835), .B($abc$9276$new_n839), .X($abc$9276$new_n843)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9775 (
        .A($abc$9276$new_n842), .B($abc$9276$new_n843), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8899)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9776 (
        .A(CPU.cli), .B($abc$9276$new_n752), .Y($abc$9276$new_n845)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9777 (
        .A($abc$9276$new_n763), .B($abc$9276$new_n779), .X($abc$9276$new_n846)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9778 (
        .A($abc$9276$new_n830), .B($abc$9276$new_n846), .X($abc$9276$new_n847)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9779 (
        .A($abc$9276$new_n845), .B($abc$9276$new_n847), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8901)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9780 (
        .A(CPU.sei), .B($abc$9276$new_n752), .Y($abc$9276$new_n849)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9781 (
        .A($abc$9276$new_n835), .B($abc$9276$new_n846), .X($abc$9276$new_n850)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9782 (
        .A($abc$9276$new_n849), .B($abc$9276$new_n850), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8903)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9783 (
        .A(CPU.clv), .B($abc$9276$new_n752), .Y($abc$9276$new_n852)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9784 (
        .A($abc$9276$new_n769), .B($abc$9276$new_n789), .X($abc$9276$new_n853)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9785 (
        .A($abc$9276$new_n853), .Y($abc$9276$new_n854)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9786 (
        .A($abc$9276$new_n835), .B($abc$9276$new_n853), .X($abc$9276$new_n855)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9787 (
        .A($abc$9276$new_n852), .B($abc$9276$new_n855), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8905)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9788 (
        .A(CPU.bit_ins), .B($abc$9276$new_n752), .Y($abc$9276$new_n857)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9789 (
        .A($abc$9276$new_n802), .B($abc$9276$new_n813), .X($abc$9276$new_n858)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9790 (
        .A($abc$9276$new_n803), .B($abc$9276$new_n813), .X($abc$9276$new_n859)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9791 (
        .A($abc$9276$new_n790), .B($abc$9276$new_n859), .X($abc$9276$new_n860)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9792 (
        .A($abc$9276$new_n752), .B($abc$9276$new_n860), .X($abc$9276$new_n861)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9793 (
        .A($abc$9276$new_n857), .B($abc$9276$new_n861), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8907)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9794 (
        .A(CPU.rotate), .B($abc$9276$new_n752), .Y($abc$9276$new_n863)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9795 (
        .A($abc$9276$new_n795), .B($abc$9276$new_n802), .X($abc$9276$new_n864)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9796 (
        .A($abc$9276$new_n815), .B($abc$9276$new_n864), .X($abc$9276$new_n865)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9797 (
        .A($abc$9276$new_n813), .B($abc$9276$new_n864), .X($abc$9276$new_n866)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9798 (
        .A($abc$9276$new_n865), .B($abc$9276$new_n866), .Y($abc$9276$new_n867)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9799 (
        .A($abc$9276$new_n752), .B($abc$9276$new_n779), .X($abc$9276$new_n868)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9800 (
        .A($abc$9276$new_n868), .Y($abc$9276$new_n869)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9801 (
        .A($abc$9276$new_n867), .B($abc$9276$new_n869), .Y($abc$9276$new_n870)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9802 (
        .A($abc$9276$new_n828), .B($abc$9276$new_n870), .X($abc$9276$new_n871)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9803 (
        .A($abc$9276$new_n779), .B($abc$9276$new_n865), .X($abc$9276$new_n872)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9804 (
        .A($abc$9276$new_n863), .B($abc$9276$new_n871), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8909)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9805 (
        .A($abc$9276$new_n846), .B($abc$9276$new_n864), .X($abc$9276$new_n874)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9806 (
        .A($abc$9276$new_n752), .B($abc$9276$new_n874), .X($abc$9276$new_n875)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9807 (
        .A(CPU.shift_right), .B($abc$9276$new_n752), .Y($abc$9276$new_n876)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9808 (
        .A($abc$9276$new_n875), .B($abc$9276$new_n876), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8911)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9809 (
        .A($abc$9276$new_n776), .B($abc$9276$new_n808), .Y($abc$9276$new_n878)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9810 (
        .A($abc$9276$new_n878), .Y($abc$9276$new_n879)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9811 (
        .A($abc$9276$new_n859), .B($abc$9276$new_n879), .X($abc$9276$new_n880)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9812 (
        .A($abc$9276$new_n880), .Y($abc$9276$new_n881)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9813 (
        .A($abc$9276$new_n769), .B($abc$9276$new_n777), .X($abc$9276$new_n882)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9814 (
        .A($abc$9276$new_n763), .B($abc$9276$new_n882), .X($abc$9276$new_n883)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9815 (
        .A($abc$9276$new_n880), .B($abc$9276$new_n883), .X($abc$9276$new_n884)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9816 (
        .A($abc$9276$new_n803), .B($abc$9276$new_n839), .X($abc$9276$new_n885)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9817 (
        .A($abc$9276$new_n775), .B($abc$9276$new_n878), .X($abc$9276$new_n886)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9818 (
        .A($abc$9276$new_n885), .B($abc$9276$new_n886), .X($abc$9276$new_n887)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9819 (
        .A($abc$9276$new_n884), .B($abc$9276$new_n887), .Y($abc$9276$new_n888)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9820 (
        .A($abc$9276$new_n795), .B($abc$9276$new_n801), .Y($abc$9276$new_n889)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9821 (
        .A($abc$9276$new_n764), .B($abc$9276$new_n786), .Y($abc$9276$new_n890)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9822 (
        .A($abc$9276$new_n889), .B($abc$9276$new_n890), .X($abc$9276$new_n891)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9823 (
        .A($abc$9276$new_n780), .B($abc$9276$new_n891), .X($abc$9276$new_n892)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9824 (
        .A($abc$9276$new_n753), .B($abc$9276$new_n892), .Y($abc$9276$new_n893)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9825 (
        .A($abc$9276$new_n888), .B($abc$9276$new_n893), .X($abc$9276$new_n894)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9826 (
        .A($abc$9276$new_n358), .B($abc$9276$new_n752), .Y($abc$9276$new_n895)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9827 (
        .A($abc$9276$new_n894), .B($abc$9276$new_n895), .Y($abc$9276$new_n896)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9828 (
        .A($abc$9276$new_n896), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8913)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9829 (
        .A(CPU.shift), .B($abc$9276$new_n752), .Y($abc$9276$new_n898)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9830 (
        .A($abc$9276$new_n870), .B($abc$9276$new_n898), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8915)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9831 (
        .A($abc$9276$new_n397), .B($abc$9276$new_n428), .Y($abc$9276$new_n900)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9832 (
        .A(in_35), .B($abc$9276$new_n900), .Y($abc$9276$new_n901)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9833 (
        .A(CPU.adc_sbc), .B($abc$9276$new_n901), .Y($abc$9276$new_n902)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9834 (
        .A($abc$9276$new_n789), .B($abc$9276$new_n827), .Y($abc$9276$new_n903)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9835 (
        .A($abc$9276$new_n889), .B($abc$9276$new_n901), .X($abc$9276$new_n904)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9836 (
        .A($abc$9276$new_n903), .B($abc$9276$new_n904), .X($abc$9276$new_n905)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9837 (
        .A($abc$9276$new_n902), .B($abc$9276$new_n905), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8917)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9838 (
        .A(CPU.adc_bcd), .B($abc$9276$new_n901), .Y($abc$9276$new_n907)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9839 (
        .A(CPU.D), .B($abc$9276$new_n780), .Y($abc$9276$new_n908)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9840 (
        .A($abc$9276$new_n905), .B($abc$9276$new_n908), .X($abc$9276$new_n909)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9841 (
        .A($abc$9276$new_n907), .B($abc$9276$new_n909), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8921)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9842 (
        .A($abc$9276$new_n839), .B($abc$9276$new_n866), .X($abc$9276$new_n911)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9843 (
        .A($abc$9276$new_n828), .B($abc$9276$new_n911), .X($abc$9276$new_n912)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9844 (
        .A($abc$9276$new_n816), .B($abc$9276$new_n883), .X($abc$9276$new_n913)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9845 (
        .A($abc$9276$new_n912), .B($abc$9276$new_n913), .Y($abc$9276$new_n914)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9846 (
        .A($abc$9276$new_n753), .B($abc$9276$new_n914), .Y($abc$9276$new_n915)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9847 (
        .A(CPU.inc), .B($abc$9276$new_n752), .Y($abc$9276$new_n916)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9848 (
        .A($abc$9276$new_n915), .B($abc$9276$new_n916), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8923)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9849 (
        .A($abc$9276$new_n786), .B($abc$9276$new_n853), .X($abc$9276$new_n918)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9850 (
        .A($abc$9276$new_n752), .B($abc$9276$new_n918), .X($abc$9276$new_n919)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9851 (
        .A(CPU.load_only), .B($abc$9276$new_n752), .Y($abc$9276$new_n920)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9852 (
        .A($abc$9276$new_n919), .B($abc$9276$new_n920), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8925)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9853 (
        .A(CPU.write_back), .B($abc$9276$new_n752), .Y($abc$9276$new_n922)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9854 (
        .A($abc$9276$new_n753), .B($abc$9276$new_n853), .Y($abc$9276$new_n923)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9855 (
        .A($abc$9276$new_n866), .B($abc$9276$new_n923), .X($abc$9276$new_n924)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9856 (
        .A($abc$9276$new_n922), .B($abc$9276$new_n924), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8927)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9857 (
        .A($abc$9276$new_n858), .B($abc$9276$new_n889), .Y($abc$9276$new_n926)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9858 (
        .A(CPU.store), .B($abc$9276$new_n752), .Y($abc$9276$new_n927)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9859 (
        .A($abc$9276$new_n854), .B($abc$9276$new_n926), .Y($abc$9276$new_n928)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9860 (
        .A($abc$9276$new_n752), .B($abc$9276$new_n827), .X($abc$9276$new_n929)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9861 (
        .A($abc$9276$new_n928), .B($abc$9276$new_n929), .X($abc$9276$new_n930)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9862 (
        .A($abc$9276$new_n927), .B($abc$9276$new_n930), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8929)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9863 (
        .A($abc$9276$new_n813), .B($abc$9276$new_n879), .Y($abc$9276$new_n932)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9864 (
        .A($abc$9276$new_n889), .B($abc$9276$new_n932), .X($abc$9276$new_n933)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9865 (
        .A($abc$9276$new_n778), .B($abc$9276$new_n933), .X($abc$9276$new_n934)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9866 (
        .A($abc$9276$new_n815), .B($abc$9276$new_n889), .X($abc$9276$new_n935)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9867 (
        .A($abc$9276$new_n753), .B($abc$9276$new_n935), .Y($abc$9276$new_n936)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9868 (
        .A($abc$9276$new_n853), .B($abc$9276$new_n864), .X($abc$9276$new_n937)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9869 (
        .A($abc$9276$new_n937), .Y($abc$9276$new_n938)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9870 (
        .A($abc$9276$new_n774), .B($abc$9276$new_n853), .X($abc$9276$new_n939)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9871 (
        .A($abc$9276$new_n866), .B($abc$9276$new_n939), .X($abc$9276$new_n940)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9872 (
        .A($abc$9276$new_n934), .B($abc$9276$new_n940), .Y($abc$9276$new_n941)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9873 (
        .A($abc$9276$new_n936), .B($abc$9276$new_n941), .X($abc$9276$new_n942)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9874 (
        .A(CPU.index_y), .B($abc$9276$new_n753), .X($abc$9276$new_n943)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9875 (
        .A($abc$9276$new_n942), .B($abc$9276$new_n943), .Y($abc$9276$new_n944)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9876 (
        .A($abc$9276$new_n944), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8931)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9877 (
        .A(CPU.load_reg), .B($abc$9276$new_n753), .X($abc$9276$new_n946)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9878 (
        .A($abc$9276$new_n816), .B($abc$9276$new_n872), .Y($abc$9276$new_n947)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9879 (
        .A($abc$9276$new_n778), .B($abc$9276$new_n947), .Y($abc$9276$new_n948)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9880 (
        .A($abc$9276$new_n948), .Y($abc$9276$new_n949)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9881 (
        .A($abc$9276$new_n858), .B($abc$9276$new_n865), .Y($abc$9276$new_n950)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9882 (
        .A($abc$9276$new_n774), .B($abc$9276$new_n918), .X($abc$9276$new_n951)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9883 (
        .A($abc$9276$new_n801), .B($abc$9276$new_n853), .X($abc$9276$new_n952)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9884 (
        .A($abc$9276$new_n808), .B($abc$9276$new_n827), .X($abc$9276$new_n953)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9885 (
        .A($abc$9276$new_n814), .B($abc$9276$new_n953), .X($abc$9276$new_n954)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9886 (
        .A($abc$9276$new_n770), .B($abc$9276$new_n786), .Y($abc$9276$new_n955)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9887 (
        .A($abc$9276$new_n955), .Y($abc$9276$new_n956)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9888 (
        .A($abc$9276$new_n777), .B($abc$9276$new_n955), .X($abc$9276$new_n957)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9889 (
        .A($abc$9276$new_n882), .B($abc$9276$new_n890), .X($abc$9276$new_n958)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9890 (
        .A($abc$9276$new_n865), .B($abc$9276$new_n958), .X($abc$9276$new_n959)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9891 (
        .A($abc$9276$new_n959), .Y($abc$9276$new_n960)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9892 (
        .A($abc$9276$new_n889), .B($abc$9276$new_n956), .X($abc$9276$new_n961)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9893 (
        .A($abc$9276$new_n951), .B($abc$9276$new_n959), .Y($abc$9276$new_n962)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9894 (
        .A($abc$9276$new_n950), .B($abc$9276$new_n962), .Y($abc$9276$new_n963)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9895 (
        .A($abc$9276$new_n853), .B($abc$9276$new_n954), .X($abc$9276$new_n964)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9896 (
        .A($abc$9276$new_n802), .B($abc$9276$new_n964), .X($abc$9276$new_n965)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9897 (
        .A($abc$9276$new_n961), .B($abc$9276$new_n965), .Y($abc$9276$new_n966)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9898 (
        .A($abc$9276$new_n966), .Y($abc$9276$new_n967)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9899 (
        .A($abc$9276$new_n963), .B($abc$9276$new_n967), .Y($abc$9276$new_n968)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9900 (
        .A($abc$9276$new_n787), .B($abc$9276$new_n952), .X($abc$9276$new_n969)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9901 (
        .A($abc$9276$new_n753), .B($abc$9276$new_n969), .Y($abc$9276$new_n970)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9902 (
        .A($abc$9276$new_n968), .B($abc$9276$new_n970), .X($abc$9276$new_n971)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9903 (
        .A($abc$9276$new_n949), .B($abc$9276$new_n971), .X($abc$9276$new_n972)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9904 (
        .A($abc$9276$new_n946), .B($abc$9276$new_n972), .Y($abc$9276$new_n973)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9905 (
        .A($abc$9276$new_n973), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8933)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9906 (
        .A($abc$9276$new_n428), .B($abc$9276$new_n760), .X($abc$9276$new_n975)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9907 (
        .A($abc$9276$new_n382), .B($abc$9276$new_n400), .X($abc$9276$new_n976)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9908 (
        .A($abc$9276$new_n393), .B($abc$9276$new_n976), .X($abc$9276$new_n977)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9909 (
        .A($abc$9276$new_n977), .Y($abc$9276$new_n978)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9910 (
        .A(CPU.backwards), .B(CPU.ALU.CO), .X($abc$9276$new_n979)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9911 (
        .A(CPU.backwards), .B(CPU.ALU.CO), .Y($abc$9276$new_n980)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9912 (
        .A($abc$9276$new_n979), .B($abc$9276$new_n980), .Y($abc$9276$new_n981)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9913 (
        .A($abc$9276$new_n978), .B($abc$9276$new_n981), .Y($abc$9276$new_n982)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9914 (
        .A($abc$9276$new_n975), .B($abc$9276$new_n982), .Y($abc$9276$new_n983)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9915 (
        .A($abc$9276$new_n410), .B($abc$9276$new_n736), .Y($abc$9276$new_n984)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9916 (
        .A($abc$9276$new_n393), .B($abc$9276$new_n728), .X($abc$9276$new_n985)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9917 (
        .A($abc$9276$new_n985), .Y($abc$9276$new_n986)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9918 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n735), .X($abc$9276$new_n987)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9919 (
        .A($abc$9276$new_n985), .B($abc$9276$new_n987), .Y($abc$9276$new_n988)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9920 (
        .A($abc$9276$new_n984), .B($abc$9276$new_n988), .X($abc$9276$new_n989)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9921 (
        .A($abc$9276$new_n983), .B($abc$9276$new_n989), .X($abc$9276$new_n990)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9922 (
        .A(oeb_0), .B($abc$9276$new_n977), .Y($abc$9276$new_n991)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9923 (
        .A($abc$9276$new_n429), .B($abc$9276$new_n991), .X($abc$9276$new_n992)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9924 (
        .A($abc$9276$new_n992), .Y($abc$9276$new_n993)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9925 (
        .A($abc$9276$new_n388), .B($abc$9276$new_n728), .X($abc$9276$new_n994)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9926 (
        .A($abc$9276$new_n386), .B($abc$9276$new_n399), .X($abc$9276$new_n995)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9927 (
        .A($abc$9276$new_n380), .B($abc$9276$new_n995), .X($abc$9276$new_n996)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9928 (
        .A($abc$9276$new_n994), .B($abc$9276$new_n996), .Y($abc$9276$new_n997)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9929 (
        .A($abc$9276$new_n388), .B($abc$9276$new_n995), .X($abc$9276$new_n998)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9930 (
        .A($abc$9276$new_n998), .Y($abc$9276$new_n999)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9931 (
        .A($abc$9276$new_n997), .B($abc$9276$new_n999), .X($abc$9276$new_n1000)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9932 (
        .A($abc$9276$new_n393), .B($abc$9276$new_n401), .X($abc$9276$new_n1001)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9933 (
        .A($abc$9276$new_n1001), .Y($abc$9276$new_n1002)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9934 (
        .A($abc$9276$new_n384), .B($abc$9276$new_n431), .Y($abc$9276$new_n1003)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9935 (
        .A($abc$9276$new_n394), .B($abc$9276$new_n1003), .Y($abc$9276$new_n1004)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9936 (
        .A($abc$9276$new_n1001), .B($abc$9276$new_n1004), .Y($abc$9276$new_n1005)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9937 (
        .A($abc$9276$new_n1000), .B($abc$9276$new_n1005), .X($abc$9276$new_n1006)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9938 (
        .A($abc$9276$new_n993), .B($abc$9276$new_n1006), .X($abc$9276$new_n1007)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9939 (
        .A($abc$9276$new_n990), .B($abc$9276$new_n1007), .X($abc$9276$new_n1008)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9940 (
        .A($abc$9276$new_n388), .B($abc$9276$new_n735), .X($abc$9276$new_n1009)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9941 (
        .A($abc$9276$new_n987), .B($abc$9276$new_n1009), .Y($abc$9276$new_n1010)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9942 (
        .A($abc$9276$new_n1000), .B($abc$9276$new_n1010), .X($abc$9276$new_n1011)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9943 (
        .A($abc$9276$new_n387), .B($abc$9276$new_n393), .X($abc$9276$new_n1012)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9944 (
        .A($abc$9276$new_n1012), .Y($abc$9276$new_n1013)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9945 (
        .A($abc$9276$new_n428), .B($abc$9276$new_n977), .Y($abc$9276$new_n1014)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9946 (
        .A($abc$9276$new_n1013), .B($abc$9276$new_n1014), .X($abc$9276$new_n1015)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9947 (
        .A($abc$9276$new_n986), .B($abc$9276$new_n1015), .X($abc$9276$new_n1016)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9948 (
        .A($abc$9276$new_n1011), .B($abc$9276$new_n1016), .X($abc$9276$new_n1017)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9949 (
        .A($abc$9276$new_n975), .B($abc$9276$new_n1017), .Y($abc$9276$new_n1018)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9950 (
        .A($abc$9276$new_n986), .B($abc$9276$new_n1018), .X($abc$9276$new_n1019)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9951 (
        .A(CPU.PC), .B($abc$9276$new_n1019), .Y($abc$9276$new_n1020)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9952 (
        .A(CPU.ADD), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1021)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9953 (
        .A($abc$9276$new_n428), .B($abc$9276$new_n759), .X($abc$9276$new_n1022)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9954 (
        .A($abc$9276$new_n1022), .Y($abc$9276$new_n1023)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9955 (
        .A(CPU.ABL), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1024)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9956 (
        .A($abc$9276$new_n373), .B($abc$9276$new_n977), .X($abc$9276$new_n1025)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9957 (
        .A($abc$9276$new_n1024), .B($abc$9276$new_n1025), .Y($abc$9276$new_n1026)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9958 (
        .A($abc$9276$new_n1026), .Y($abc$9276$new_n1027)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9959 (
        .A($abc$9276$new_n1021), .B($abc$9276$new_n1027), .Y($abc$9276$new_n1028)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9960 (
        .A($abc$9276$new_n1028), .Y($abc$9276$new_n1029)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9961 (
        .A($abc$9276$new_n1020), .B($abc$9276$new_n1029), .Y($abc$9276$new_n1030)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9962 (
        .A($abc$9276$new_n1008), .B($abc$9276$new_n1030), .Y($abc$9276$new_n1031)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9963 (
        .A($abc$9276$new_n1031), .Y($abc$9276$new_n1032)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9964 (
        .A($abc$9276$new_n1008), .B($abc$9276$new_n1030), .X($abc$9276$new_n1033)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9965 (
        .A($abc$9276$new_n1031), .B($abc$9276$new_n1033), .Y($abc$9276$new_n1034)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9966 (
        .A(in_35), .B($abc$9276$new_n1034), .Y($abc$9276$new_n1035)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9967 (
        .A(CPU.PC), .B(in_35), .X($abc$9276$new_n1036)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9968 (
        .A($abc$9276$new_n1035), .B($abc$9276$new_n1036), .Y($abc$9276$new_n1037)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9969 (
        .A($abc$9276$new_n1037), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8935)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9970 (
        .A(CPU.PC), .B($abc$9276$new_n1019), .Y($abc$9276$new_n1039)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9971 (
        .A(CPU.ADD), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1040)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9972 (
        .A(CPU.ABL), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1041)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9973 (
        .A(CPU.ADD), .B($abc$9276$new_n978), .Y($abc$9276$new_n1042)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9974 (
        .A($abc$9276$new_n1042), .Y($abc$9276$new_n1043)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9975 (
        .A($flatten\CPU.$procmux$715.B), .B($abc$9276$new_n1013), .Y($abc$9276$new_n1044)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9976 (
        .A($abc$9276$new_n1041), .B($abc$9276$new_n1044), .Y($abc$9276$new_n1045)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9977 (
        .A($abc$9276$new_n1040), .B($abc$9276$new_n1042), .Y($abc$9276$new_n1046)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9978 (
        .A($abc$9276$new_n1045), .B($abc$9276$new_n1046), .X($abc$9276$new_n1047)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9979 (
        .A($abc$9276$new_n1047), .Y($abc$9276$new_n1048)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9980 (
        .A($abc$9276$new_n1039), .B($abc$9276$new_n1048), .Y($abc$9276$new_n1049)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9981 (
        .A($abc$9276$new_n1032), .B($abc$9276$new_n1049), .Y($abc$9276$new_n1050)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9982 (
        .A($abc$9276$new_n1050), .Y($abc$9276$new_n1051)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9983 (
        .A($abc$9276$new_n1032), .B($abc$9276$new_n1049), .X($abc$9276$new_n1052)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9984 (
        .A($abc$9276$new_n1050), .B($abc$9276$new_n1052), .Y($abc$9276$new_n1053)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9985 (
        .A(in_35), .B($abc$9276$new_n1053), .Y($abc$9276$new_n1054)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9986 (
        .A(in_35), .B(CPU.PC), .X($abc$9276$new_n1055)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9987 (
        .A($abc$9276$new_n1054), .B($abc$9276$new_n1055), .Y($abc$9276$new_n1056)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9988 (
        .A($abc$9276$new_n1056), .Y($abc$9276$auto$rtlil.cc:3205:MuxGate$8937)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9989 (
        .A(CPU.PC), .B($abc$9276$new_n1019), .Y($abc$9276$new_n1058)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9990 (
        .A(CPU.ADD), .B($abc$9276$new_n1011), .Y($abc$9276$new_n1059)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9991 (
        .A($abc$9276$new_n1059), .Y($abc$9276$new_n1060)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9992 (
        .A(CPU.ABL), .B($abc$9276$new_n1023), .Y($abc$9276$new_n1061)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9993 (
        .A($abc$9276$new_n374), .B($abc$9276$new_n977), .X($abc$9276$new_n1062)
    );

    sky130_fd_sc_hd__clkinv_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9994 (
        .A($abc$9276$new_n1062), .Y($abc$9276$new_n1063)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9995 (
        .A($abc$9276$new_n351), .B(CPU.res), .Y($abc$9276$new_n1064)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9996 (
        .A(CPU.res), .B($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9264), .X($abc$9276$new_n1065)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9997 (
        .A($abc$9276$new_n1064), .B($abc$9276$new_n1065), .Y($abc$9276$new_n1066)
    );

    sky130_fd_sc_hd__or2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9998 (
        .A($abc$9276$new_n1012), .B($abc$9276$new_n1066), .X($abc$9276$new_n1067)
    );

    sky130_fd_sc_hd__nand2_2 $abc$9276$auto$blifparse.cc:396:parse_blif$9999 (
        .A($abc$9276$new_n1061), .B($abc$9276$new_n1067), .Y($abc$9276$new_n1068)
    );

    sky130_fd_sc_hd__conb_1 $auto$hilomap.cc:40:hilomap_worker$12031 (
        .HI($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__conb_1 $auto$hilomap.cc:40:hilomap_worker$8815 (
        .HI(oeb_16)
    );

    sky130_fd_sc_hd__conb_1 $auto$hilomap.cc:48:hilomap_worker$8817 (
        .LO(oeb_0)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11708 (
        .A(CPU.Z), .Y($flatten\CPU.$procmux$291.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11709 (
        .A(CPU.C), .Y($flatten\CPU.$procmux$291.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11710 (
        .A(CPU.V), .Y($flatten\CPU.$procmux$291.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11711 (
        .A(CPU.N), .Y($flatten\CPU.$procmux$291.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11712 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11713 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11714 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11715 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11716 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11717 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11718 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11719 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11720 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11721 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11722 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11723 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11724 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11725 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11726 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11727 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11728 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11729 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11730 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11731 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11732 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11733 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11734 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11735 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11736 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11737 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11738 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11739 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11740 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11741 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11742 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11743 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11744 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11745 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11746 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11747 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11748 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11749 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11750 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11751 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11752 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11753 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11754 (
        .A($flatten\CPU.$procmux$415.B), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11755 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11756 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11757 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11758 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11759 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11760 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11761 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11762 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11763 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11764 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11765 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11766 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11767 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11768 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11769 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11770 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11771 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11772 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11773 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11774 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11775 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11776 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11777 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11778 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11779 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11780 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11781 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11782 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11783 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11784 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11785 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11786 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11787 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11788 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11789 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11790 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11791 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11792 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11793 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11794 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11795 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11796 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11797 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11798 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11799 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11800 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11801 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11802 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11803 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11804 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11805 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11806 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11807 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11808 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11809 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11810 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11811 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11812 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11813 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11814 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11815 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11816 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11817 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11818 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11819 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11820 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11821 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11822 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11823 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11824 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11825 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11826 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11827 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11828 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11829 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11830 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11831 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11832 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11833 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11834 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11835 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11836 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11837 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11838 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11839 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11840 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11841 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11842 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11843 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11844 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11845 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11846 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11847 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11848 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11849 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11850 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11851 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11852 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11853 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11854 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11855 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11856 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11857 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11858 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11859 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11860 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11861 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11862 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11863 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11864 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11865 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11866 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11867 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11868 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11869 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11870 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11871 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11872 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11873 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11874 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11875 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11876 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11877 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11878 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11879 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11880 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11881 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11882 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11883 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11884 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11885 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11886 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11887 (
        .A(CPU.write_back), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11888 (
        .A($flatten\CPU.$procmux$415.B), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11889 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11890 (
        .A(CPU.write_back), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11891 (
        .A($flatten\CPU.$procmux$415.B), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11892 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11893 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11894 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11895 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11896 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11897 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11898 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11899 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11900 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11901 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11902 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11903 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11904 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11905 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11906 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11907 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11908 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11909 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11910 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11911 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11912 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11913 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$415.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11914 (
        .A(oeb_0), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11915 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11916 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11917 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11918 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11919 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11920 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11921 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11922 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11923 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11924 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11925 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11926 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11927 (
        .A(oeb_16), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11928 (
        .A(CPU.PC), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11929 (
        .A(CPU.PC), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11930 (
        .A(CPU.PC), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11931 (
        .A(CPU.PC), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11932 (
        .A(CPU.PC), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11933 (
        .A(CPU.PC), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11934 (
        .A(CPU.PC), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11935 (
        .A(CPU.PC), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11936 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11937 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11938 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11939 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11940 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11941 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11942 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11943 (
        .A(CPU.ALU.N), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11944 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11945 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11946 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11947 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11948 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11949 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11950 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11951 (
        .A(CPU.ALU.N), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11952 (
        .A(CPU.ABH), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11953 (
        .A(CPU.ABH), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11954 (
        .A(CPU.ABH), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11955 (
        .A(CPU.ABH), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11956 (
        .A(CPU.ABH), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11957 (
        .A(CPU.ABH), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11958 (
        .A(CPU.ABH), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11959 (
        .A(CPU.ABH), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11960 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11961 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11962 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11963 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11964 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11965 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11966 (
        .A(CPU.ADD), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11967 (
        .A(CPU.ALU.N), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11968 (
        .A(CPU.DIMUX), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11969 (
        .A(CPU.DIMUX), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11970 (
        .A(CPU.DIMUX), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11971 (
        .A(CPU.DIMUX), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11972 (
        .A(CPU.DIMUX), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11973 (
        .A(CPU.DIMUX), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11974 (
        .A(CPU.DIMUX), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11975 (
        .A(CPU.DIMUX), .Y($flatten\CPU.$procmux$715.B)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11976 (
        .A(CPU.ALU.N), .Y(CPU.ADD)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11977 (
        .A(oeb_0), .Y(oeb_1)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11978 (
        .A(oeb_0), .Y(oeb_10)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11979 (
        .A(oeb_0), .Y(oeb_11)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11980 (
        .A(oeb_0), .Y(oeb_12)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11981 (
        .A(oeb_0), .Y(oeb_13)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11982 (
        .A(oeb_0), .Y(oeb_14)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11983 (
        .A(oeb_0), .Y(oeb_15)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11984 (
        .A(oeb_16), .Y(oeb_17)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11985 (
        .A(oeb_16), .Y(oeb_18)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11986 (
        .A(oeb_16), .Y(oeb_19)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11987 (
        .A(oeb_0), .Y(oeb_2)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11988 (
        .A(oeb_16), .Y(oeb_20)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11989 (
        .A(oeb_16), .Y(oeb_21)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11990 (
        .A(oeb_16), .Y(oeb_22)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11991 (
        .A(oeb_16), .Y(oeb_23)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11992 (
        .A(oeb_0), .Y(oeb_24)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11993 (
        .A(oeb_0), .Y(oeb_25)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11994 (
        .A(oeb_0), .Y(oeb_26)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11995 (
        .A(oeb_0), .Y(oeb_27)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11996 (
        .A(oeb_0), .Y(oeb_28)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11997 (
        .A(oeb_0), .Y(oeb_29)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11998 (
        .A(oeb_0), .Y(oeb_3)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$11999 (
        .A(oeb_0), .Y(oeb_30)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12000 (
        .A(oeb_0), .Y(oeb_31)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12001 (
        .A(oeb_0), .Y(oeb_32)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12002 (
        .A(oeb_16), .Y(oeb_33)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12003 (
        .A(oeb_16), .Y(oeb_34)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12004 (
        .A(oeb_16), .Y(oeb_35)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12005 (
        .A(oeb_16), .Y(oeb_36)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12006 (
        .A(oeb_16), .Y(oeb_37)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12007 (
        .A(oeb_16), .Y(oeb_38)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12008 (
        .A(oeb_16), .Y(oeb_39)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12009 (
        .A(oeb_0), .Y(oeb_4)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12010 (
        .A(oeb_0), .Y(oeb_5)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12011 (
        .A(oeb_0), .Y(oeb_6)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12012 (
        .A(oeb_0), .Y(oeb_7)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12013 (
        .A(oeb_0), .Y(oeb_8)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12014 (
        .A(oeb_0), .Y(oeb_9)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12015 (
        .A(oeb_0), .Y(out_16)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12016 (
        .A(oeb_0), .Y(out_17)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12017 (
        .A(oeb_0), .Y(out_18)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12018 (
        .A(oeb_0), .Y(out_19)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12019 (
        .A(oeb_0), .Y(out_20)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12020 (
        .A(oeb_0), .Y(out_21)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12021 (
        .A(oeb_0), .Y(out_22)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12022 (
        .A(oeb_0), .Y(out_23)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12023 (
        .A(oeb_0), .Y(out_33)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12024 (
        .A(oeb_0), .Y(out_34)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12025 (
        .A(oeb_0), .Y(out_35)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12026 (
        .A(oeb_0), .Y(out_36)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12027 (
        .A(oeb_0), .Y(out_37)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12028 (
        .A(oeb_0), .Y(out_38)
    );

    sky130_fd_sc_hd__clkbuf_4 $auto$insbuf.cc:97:execute$12029 (
        .A(oeb_0), .Y(out_39)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4105 (
        .CLK(cts_net_3140), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8819), .Q(CPU.AXYS[3]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9263), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4106 (
        .CLK(cts_net_3144), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8821), .Q(CPU.AXYS[3]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9262), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4107 (
        .CLK(cts_net_3159), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8823), .Q(CPU.AXYS[3]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9261), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4108 (
        .CLK(cts_net_3186), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8825), .Q(CPU.AXYS[3]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9260), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4109 (
        .CLK(cts_net_3156), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8827), .Q(CPU.AXYS[3]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9259), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4110 (
        .CLK(cts_net_3141), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8829), .Q(CPU.AXYS[3]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9258), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4111 (
        .CLK(cts_net_3182), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8831), .Q(CPU.AXYS[3]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9257), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4112 (
        .CLK(cts_net_3128), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8833), .Q(CPU.AXYS[3]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9256), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4907 (
        .CLK(cts_net_3158), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8835), .Q(CPU.AXYS[2]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9255), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4908 (
        .CLK(cts_net_3141), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8837), .Q(CPU.AXYS[2]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9254), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4909 (
        .CLK(cts_net_3166), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8839), .Q(CPU.AXYS[2]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9253), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4910 (
        .CLK(cts_net_3121), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8841), .Q(CPU.AXYS[2]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9252), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4911 (
        .CLK(cts_net_3167), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8843), .Q(CPU.AXYS[2]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9251), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4912 (
        .CLK(cts_net_3159), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8845), .Q(CPU.AXYS[2]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9250), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4913 (
        .CLK(cts_net_3129), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8847), .Q(CPU.AXYS[2]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9249), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4914 (
        .CLK(cts_net_3124), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8849), .Q(CPU.AXYS[2]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9248), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4931 (
        .CLK(cts_net_3131), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8851), .Q(CPU.AXYS[1]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9247), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4932 (
        .CLK(cts_net_3131), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8853), .Q(CPU.AXYS[1]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9246), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4933 (
        .CLK(cts_net_3140), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8855), .Q(CPU.AXYS[1]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9245), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4934 (
        .CLK(cts_net_3167), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8857), .Q(CPU.AXYS[1]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9244), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4935 (
        .CLK(cts_net_3144), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8859), .Q(CPU.AXYS[1]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9243), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4936 (
        .CLK(cts_net_3155), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8861), .Q(CPU.AXYS[1]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9242), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4937 (
        .CLK(cts_net_3155), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8863), .Q(CPU.AXYS[1]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9241), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4938 (
        .CLK(cts_net_3144), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8865), .Q(CPU.AXYS[1]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9240), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4979 (
        .CLK(cts_net_3145), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8867), .Q(CPU.AXYS[0]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9239), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4980 (
        .CLK(cts_net_3132), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8869), .Q(CPU.AXYS[0]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9238), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4981 (
        .CLK(cts_net_3128), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8871), .Q(CPU.AXYS[0]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9237), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4982 (
        .CLK(cts_net_3145), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8873), .Q(CPU.AXYS[0]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9236), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4983 (
        .CLK(cts_net_3138), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8875), .Q(CPU.AXYS[0]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9235), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4984 (
        .CLK(cts_net_3185), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8877), .Q(CPU.AXYS[0]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9234), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4985 (
        .CLK(cts_net_3182), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8879), .Q(CPU.AXYS[0]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9233), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$4986 (
        .CLK(cts_net_3148), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8881), .Q(CPU.AXYS[0]), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9232), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5134 (
        .CLK(cts_net_3190), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8883), .Q(CPU.V), .Q_N($flatten\CPU.$procmux$291.B), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5135 (
        .CLK(cts_net_3174), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8887), .Q(CPU.NMI_edge), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9264), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5136 (
        .CLK(cts_net_3202), .D(in_34), .Q(CPU.NMI_1), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9228), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5137 (
        .CLK(cts_net_3141), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8889), .Q(CPU.plp), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9226), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5138 (
        .CLK(cts_net_3185), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8891), .Q(CPU.php), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9225), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5139 (
        .CLK(cts_net_3189), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8893), .Q(CPU.clc), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9224), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5140 (
        .CLK(cts_net_3148), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8895), .Q(CPU.sec), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9223), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5141 (
        .CLK(cts_net_3192), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8897), .Q(CPU.cld), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9222), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5142 (
        .CLK(cts_net_3147), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8899), .Q(CPU.sed), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9221), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5143 (
        .CLK(cts_net_3189), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8901), .Q(CPU.cli), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9220), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5144 (
        .CLK(cts_net_3161), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8903), .Q(CPU.sei), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9219), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5145 (
        .CLK(cts_net_3161), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8905), .Q(CPU.clv), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9218), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5146 (
        .CLK(cts_net_3202), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8907), .Q(CPU.bit_ins), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9217), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5151 (
        .CLK(cts_net_3148), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8909), .Q(CPU.rotate), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9216), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5152 (
        .CLK(cts_net_3166), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8911), .Q(CPU.shift_right), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9215), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5153 (
        .CLK(cts_net_3183), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8913), .Q(CPU.compare), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9214), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5154 (
        .CLK(cts_net_3186), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8915), .Q(CPU.shift), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9213), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5155 (
        .CLK(cts_net_3167), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8917), .Q(CPU.adc_sbc), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9212), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5156 (
        .CLK(cts_net_3183), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8921), .Q(CPU.adc_bcd), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9210), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5157 (
        .CLK(cts_net_3198), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8923), .Q(CPU.inc), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9209), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5158 (
        .CLK(cts_net_3155), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8925), .Q(CPU.load_only), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9208), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5159 (
        .CLK(cts_net_3145), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8927), .Q(CPU.write_back), .Q_N($flatten\CPU.$procmux$415.B), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5160 (
        .CLK(cts_net_3192), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8929), .Q(CPU.store), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9205), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5161 (
        .CLK(cts_net_3182), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8931), .Q(CPU.index_y), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9204), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5166 (
        .CLK(cts_net_3129), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8933), .Q(CPU.load_reg), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9203), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5167 (
        .CLK(cts_net_3159), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8935), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9202), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5168 (
        .CLK(cts_net_3197), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8937), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9201), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5169 (
        .CLK(cts_net_3193), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8939), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9200), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5170 (
        .CLK(cts_net_3185), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8941), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9199), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5171 (
        .CLK(cts_net_3124), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8943), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9198), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5172 (
        .CLK(cts_net_3176), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8945), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9197), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5173 (
        .CLK(cts_net_3198), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8947), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9196), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5174 (
        .CLK(cts_net_3198), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8949), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9195), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5175 (
        .CLK(cts_net_3190), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8951), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9194), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5176 (
        .CLK(cts_net_3176), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8953), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9193), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5177 (
        .CLK(cts_net_3200), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8955), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9192), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5178 (
        .CLK(cts_net_3202), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8957), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9191), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5179 (
        .CLK(cts_net_3190), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8959), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9190), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5180 (
        .CLK(cts_net_3162), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8961), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9189), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5181 (
        .CLK(cts_net_3197), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8963), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9188), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5182 (
        .CLK(cts_net_3189), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8965), .Q(CPU.PC), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9187), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5183 (
        .CLK(cts_net_3123), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8969), .Q(CPU.res), .Q_N($flatten\CPU.$procmux$715.B), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5189 (
        .CLK(cts_net_3200), .D(CPU.DIMUX), .Q(CPU.DIHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9268), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5190 (
        .CLK(cts_net_3162), .D(CPU.DIMUX), .Q(CPU.DIHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9269), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5191 (
        .CLK(cts_net_3169), .D(CPU.DIMUX), .Q(CPU.DIHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9270), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5192 (
        .CLK(cts_net_3193), .D(CPU.DIMUX), .Q(CPU.DIHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9271), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5193 (
        .CLK(cts_net_3200), .D(CPU.DIMUX), .Q(CPU.DIHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9272), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5194 (
        .CLK(cts_net_3192), .D(CPU.DIMUX), .Q(CPU.DIHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9273), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5195 (
        .CLK(cts_net_3147), .D(CPU.DIMUX), .Q(CPU.DIHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9274), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5196 (
        .CLK(cts_net_3166), .D(CPU.DIMUX), .Q(CPU.DIHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9186), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5197 (
        .CLK(cts_net_3193), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8971), .Q(CPU.cond_code), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9184), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5198 (
        .CLK(cts_net_3202), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8973), .Q(CPU.cond_code), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9182), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5199 (
        .CLK(cts_net_3162), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8975), .Q(CPU.cond_code), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9180), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5200 (
        .CLK(cts_net_3173), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8979), .Q(CPU.IRHOLD_valid), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9179), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5201 (
        .CLK(cts_net_3124), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8981), .Q(CPU.D), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9178), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5202 (
        .CLK(cts_net_3147), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8983), .Q(CPU.N), .Q_N($flatten\CPU.$procmux$291.B), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5203 (
        .CLK(cts_net_3132), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8987), .Q(CPU.I), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9174), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5204 (
        .CLK(cts_net_3138), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8989), .Q(CPU.Z), .Q_N($flatten\CPU.$procmux$291.B), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5205 (
        .CLK(cts_net_3123), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8991), .Q(CPU.C), .Q_N($flatten\CPU.$procmux$291.B), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5206 (
        .CLK(cts_net_3162), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8993), .Q(CPU.backwards), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9169), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5207 (
        .CLK(cts_net_3183), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8995), .Q(CPU.ABL), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9168), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5208 (
        .CLK(cts_net_3131), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8997), .Q(CPU.ABL), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9167), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5209 (
        .CLK(cts_net_3186), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$8999), .Q(CPU.ABL), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9166), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5210 (
        .CLK(cts_net_3129), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9001), .Q(CPU.ABL), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9165), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5211 (
        .CLK(cts_net_3158), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9003), .Q(CPU.ABL), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9164), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5212 (
        .CLK(cts_net_3156), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9005), .Q(CPU.ABL), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9163), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5213 (
        .CLK(cts_net_3121), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9007), .Q(CPU.ABL), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9162), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5214 (
        .CLK(cts_net_3167), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9009), .Q(CPU.ABL), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9275), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5215 (
        .CLK(cts_net_3132), .D($abc$9276$flatten\CPU.$0\adj_bcd[0:0]), .Q(CPU.adj_bcd), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9160), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5216 (
        .CLK(cts_net_3150), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9011), .Q(CPU.ABH), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9159), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5217 (
        .CLK(cts_net_3137), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9013), .Q(CPU.ABH), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9158), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5218 (
        .CLK(cts_net_3151), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9015), .Q(CPU.ABH), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9157), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5219 (
        .CLK(cts_net_3151), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9017), .Q(CPU.ABH), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9156), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5220 (
        .CLK(cts_net_3120), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9019), .Q(CPU.ABH), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9155), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5221 (
        .CLK(cts_net_3150), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9021), .Q(CPU.ABH), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9154), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5222 (
        .CLK(cts_net_3151), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9023), .Q(CPU.ABH), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9153), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5223 (
        .CLK(cts_net_3125), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9025), .Q(CPU.ABH), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9152), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5224 (
        .CLK(cts_net_3176), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9027), .Q(CPU.IRHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9151), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5225 (
        .CLK(cts_net_3170), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9029), .Q(CPU.IRHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9150), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5226 (
        .CLK(cts_net_3178), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9031), .Q(CPU.IRHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9149), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5227 (
        .CLK(cts_net_3174), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9033), .Q(CPU.IRHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9148), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5228 (
        .CLK(cts_net_3201), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9035), .Q(CPU.IRHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9147), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5229 (
        .CLK(cts_net_3174), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9037), .Q(CPU.IRHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9146), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5230 (
        .CLK(cts_net_3173), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9039), .Q(CPU.IRHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9145), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5231 (
        .CLK(cts_net_3203), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9041), .Q(CPU.IRHOLD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9144), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5232 (
        .CLK(cts_net_3177), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9043), .Q(CPU.state), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9142), .RESET_B(rst_n), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5233 (
        .CLK(cts_net_3169), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9045), .Q(CPU.state), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9140), .RESET_B(rst_n), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5234 (
        .CLK(cts_net_3125), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9047), .Q(CPU.state), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9138), .RESET_B(rst_n), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5235 (
        .CLK(cts_net_3177), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9049), .Q(CPU.state), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9136), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B(rst_n)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5236 (
        .CLK(cts_net_3169), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9051), .Q(CPU.state), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9134), .RESET_B(rst_n), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$5237 (
        .CLK(cts_net_3125), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9053), .Q(CPU.state), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9132), .RESET_B(rst_n), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8804 (
        .CLK(cts_net_3174), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9057), .Q(CPU.dst_reg), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9131), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8805 (
        .CLK(cts_net_3137), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9061), .Q(CPU.dst_reg), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9130), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8806 (
        .CLK(cts_net_3121), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9065), .Q(CPU.src_reg), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9129), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8807 (
        .CLK(cts_net_3140), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9069), .Q(CPU.src_reg), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9128), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8808 (
        .CLK(cts_net_3138), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9073), .Q(CPU.op), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9127), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8809 (
        .CLK(cts_net_3170), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9077), .Q(CPU.op), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9126), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8810 (
        .CLK(cts_net_3170), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9081), .Q(CPU.op), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9125), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.$auto$ff.cc:266:slice$8811 (
        .CLK(cts_net_3151), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9085), .Q(CPU.op), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9124), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7456 (
        .CLK(cts_net_3170), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9087), .Q(CPU.ALU.BI7), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9123), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7679 (
        .CLK(cts_net_3177), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9089), .Q(CPU.ALU.N), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9122), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7680 (
        .CLK(cts_net_3177), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9091), .Q(CPU.ALU.HC), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9120), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7681 (
        .CLK(cts_net_3176), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9093), .Q(CPU.ADD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9119), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7682 (
        .CLK(cts_net_3201), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9095), .Q(CPU.ADD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9118), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7683 (
        .CLK(cts_net_3201), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9097), .Q(CPU.ADD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9117), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7684 (
        .CLK(cts_net_3203), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9099), .Q(CPU.ADD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9116), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7685 (
        .CLK(cts_net_3173), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9101), .Q(CPU.ADD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9115), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7686 (
        .CLK(cts_net_3120), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9103), .Q(CPU.ADD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9114), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7687 (
        .CLK(cts_net_3169), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9105), .Q(CPU.ADD), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9113), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7689 (
        .CLK(cts_net_3203), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9107), .Q(CPU.ALU.AI7), .Q_N($auto$dfflibmap.cc:532:dfflibmap$9112), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__dfbbp_1 $flatten\CPU.\ALU.$auto$ff.cc:266:slice$7690 (
        .CLK(cts_net_3173), .D($abc$9276$auto$rtlil.cc:3205:MuxGate$9109), .Q(CPU.ALU.CO), .Q_N($abc$9276$auto$dfflibmap.cc:532:dfflibmap$9110), .RESET_B($auto$hilomap.cc:39:hilomap_worker$12030), .SET_B($auto$hilomap.cc:39:hilomap_worker$12030)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_0_503_257 (
        .A(clk), .X(cts_net_3116)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_1_531_410 (
        .A(cts_net_3116), .X(cts_net_3117)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_2_517_440 (
        .A(cts_net_3117), .X(cts_net_3118)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_517_453 (
        .A(cts_net_3118), .X(cts_net_3119)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_461 (
        .A(cts_net_3119), .X(cts_net_3120)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_448 (
        .A(cts_net_3119), .X(cts_net_3121)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_517_426 (
        .A(cts_net_3118), .X(cts_net_3122)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_434 (
        .A(cts_net_3122), .X(cts_net_3123)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_421 (
        .A(cts_net_3122), .X(cts_net_3124)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_2_545_404 (
        .A(cts_net_3117), .X(cts_net_3125)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_2_517_383 (
        .A(cts_net_3117), .X(cts_net_3126)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_517_399 (
        .A(cts_net_3126), .X(cts_net_3127)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_407 (
        .A(cts_net_3127), .X(cts_net_3128)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_393 (
        .A(cts_net_3127), .X(cts_net_3129)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_517_369 (
        .A(cts_net_3126), .X(cts_net_3130)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_377 (
        .A(cts_net_3130), .X(cts_net_3131)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_361 (
        .A(cts_net_3130), .X(cts_net_3132)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_1_476_385 (
        .A(cts_net_3116), .X(cts_net_3133)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_2_489_448 (
        .A(cts_net_3133), .X(cts_net_3134)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_489_481 (
        .A(cts_net_3134), .X(cts_net_3135)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_489_497 (
        .A(cts_net_3135), .X(cts_net_3136)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_505 (
        .A(cts_net_3136), .X(cts_net_3137)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_491 (
        .A(cts_net_3136), .X(cts_net_3138)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_489_467 (
        .A(cts_net_3135), .X(cts_net_3139)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_475 (
        .A(cts_net_3139), .X(cts_net_3140)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_459 (
        .A(cts_net_3139), .X(cts_net_3141)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_489_418 (
        .A(cts_net_3134), .X(cts_net_3142)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_489_434 (
        .A(cts_net_3142), .X(cts_net_3143)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_442 (
        .A(cts_net_3143), .X(cts_net_3144)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_426 (
        .A(cts_net_3143), .X(cts_net_3145)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_489_402 (
        .A(cts_net_3142), .X(cts_net_3146)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_410 (
        .A(cts_net_3146), .X(cts_net_3147)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_393 (
        .A(cts_net_3146), .X(cts_net_3148)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_2_462_410 (
        .A(cts_net_3133), .X(cts_net_3149)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_462_423 (
        .A(cts_net_3149), .X(cts_net_3150)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_462_402 (
        .A(cts_net_3149), .X(cts_net_3151)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_2_489_323 (
        .A(cts_net_3133), .X(cts_net_3152)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_489_358 (
        .A(cts_net_3152), .X(cts_net_3153)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_489_372 (
        .A(cts_net_3153), .X(cts_net_3154)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_377 (
        .A(cts_net_3154), .X(cts_net_3155)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_364 (
        .A(cts_net_3154), .X(cts_net_3156)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_489_345 (
        .A(cts_net_3153), .X(cts_net_3157)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_353 (
        .A(cts_net_3157), .X(cts_net_3158)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_339 (
        .A(cts_net_3157), .X(cts_net_3159)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_489_287 (
        .A(cts_net_3152), .X(cts_net_3160)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_489_309 (
        .A(cts_net_3160), .X(cts_net_3161)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_489_271 (
        .A(cts_net_3160), .X(cts_net_3162)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_1_517_165 (
        .A(cts_net_3116), .X(cts_net_3163)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_2_517_209 (
        .A(cts_net_3163), .X(cts_net_3164)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_517_230 (
        .A(cts_net_3164), .X(cts_net_3165)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_241 (
        .A(cts_net_3165), .X(cts_net_3166)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_222 (
        .A(cts_net_3165), .X(cts_net_3167)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_517_189 (
        .A(cts_net_3164), .X(cts_net_3168)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_200 (
        .A(cts_net_3168), .X(cts_net_3169)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_179 (
        .A(cts_net_3168), .X(cts_net_3170)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_2_517_124 (
        .A(cts_net_3163), .X(cts_net_3171)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_517_146 (
        .A(cts_net_3171), .X(cts_net_3172)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_157 (
        .A(cts_net_3172), .X(cts_net_3173)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_135 (
        .A(cts_net_3172), .X(cts_net_3174)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_517_102 (
        .A(cts_net_3171), .X(cts_net_3175)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_113 (
        .A(cts_net_3175), .X(cts_net_3176)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_517_92 (
        .A(cts_net_3175), .X(cts_net_3177)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_1_476_132 (
        .A(cts_net_3116), .X(cts_net_3178)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_2_489_195 (
        .A(cts_net_3178), .X(cts_net_3179)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_489_228 (
        .A(cts_net_3179), .X(cts_net_3180)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_489_244 (
        .A(cts_net_3180), .X(cts_net_3181)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_252 (
        .A(cts_net_3181), .X(cts_net_3182)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_236 (
        .A(cts_net_3181), .X(cts_net_3183)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_489_211 (
        .A(cts_net_3180), .X(cts_net_3184)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_219 (
        .A(cts_net_3184), .X(cts_net_3185)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_203 (
        .A(cts_net_3184), .X(cts_net_3186)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_489_162 (
        .A(cts_net_3179), .X(cts_net_3187)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_489_179 (
        .A(cts_net_3187), .X(cts_net_3188)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_187 (
        .A(cts_net_3188), .X(cts_net_3189)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_170 (
        .A(cts_net_3188), .X(cts_net_3190)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_489_146 (
        .A(cts_net_3187), .X(cts_net_3191)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_154 (
        .A(cts_net_3191), .X(cts_net_3192)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_138 (
        .A(cts_net_3191), .X(cts_net_3193)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_2_489_67 (
        .A(cts_net_3178), .X(cts_net_3194)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_489_100 (
        .A(cts_net_3194), .X(cts_net_3195)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_489_116 (
        .A(cts_net_3195), .X(cts_net_3196)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_124 (
        .A(cts_net_3196), .X(cts_net_3197)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_111 (
        .A(cts_net_3196), .X(cts_net_3198)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_4_489_86 (
        .A(cts_net_3195), .X(cts_net_3199)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_94 (
        .A(cts_net_3199), .X(cts_net_3200)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_5_489_78 (
        .A(cts_net_3199), .X(cts_net_3201)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_3_489_15 (
        .A(cts_net_3194), .X(cts_net_3202)
    );

    sky130_fd_sc_hd__buf_1 cts_htree_2_462_116 (
        .A(cts_net_3178), .X(cts_net_3203)
    );

endmodule