# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
#   DISTANCE MICRONS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;
USEMINSPACING OBS OFF ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

# High density, single height
SITE unithd
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.46 BY 2.72 ;
END unithd

# High density, double height
SITE unithddbl
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell

LAYER licon
  TYPE CUT ;
END licon

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.46 0.34 ;
  OFFSET 0.23 0.17 ;

  WIDTH 0.17 ;          # LI 1
  # SPACING  0.17 ;     # LI 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.17 ;
  AREA 0.0561 ;         # LI 6
  THICKNESS 0.1 ;
  EDGECAPACITANCE 40.697E-6 ;
  CAPACITANCE CPERSQDIST 36.9866E-6 ;
  RESISTANCE RPERSQ 12.8 ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 75 ) ( 0.0125 75 ) ( 0.0225 85.125 ) ( 22.5 10200 ) ) ;
END li1

LAYER mcon
  TYPE CUT ;

  WIDTH 0.17 ;                # Mcon 1
  SPACING 0.19 ;              # Mcon 2
  ENCLOSURE BELOW 0 0 ;       # Mcon 4
  ENCLOSURE ABOVE 0.03 0.06 ; # Met1 4 / Met1 5
  RESISTANCE 9.30 ;

  ANTENNADIFFAREARATIO PWL ( ( 0 3 ) ( 0.0125 3 ) ( 0.0225 3.405 ) ( 22.5 408 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.36 ; # mA per via Iavg_max at Tj = 90oC

END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 0.34 ;
  OFFSET 0.17 ;

  WIDTH 0.14 ;                     # Met1 1
  # SPACING 0.14 ;                 # Met1 2
  # SPACING 0.28 RANGE 3.001 100 ; # Met1 3b
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.14
     WIDTH 3 0.28 ;
  AREA 0.083 ;                     # Met1 6
  THICKNESS 0.35 ;
  MINENCLOSEDAREA 0.14 ;

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  EDGECAPACITANCE 40.567E-6 ;
  CAPACITANCE CPERSQDIST 25.7784E-6 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC
  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;

  RESISTANCE RPERSQ 0.125 ;
END met1

LAYER via
  TYPE CUT ;
  WIDTH 0.15 ;                  # Via 1a
  SPACING 0.17 ;                # Via 2
  ENCLOSURE BELOW 0.055 0.085 ; # Via 4a / Via 5a
  ENCLOSURE ABOVE 0.055 0.085 ; # Met2 4 / Met2 5
  RESISTANCE 4.50 ;

  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.29 ; # mA per via Iavg_max at Tj = 90oC
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.46 ;
  OFFSET 0.23 ;

  WIDTH 0.14 ;                        # Met2 1
  # SPACING  0.14 ;                   # Met2 2
  # SPACING  0.28 RANGE 3.001 100 ;   # Met2 3b
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.14
     WIDTH 3 0.28 ;
  AREA 0.0676 ;                       # Met2 6
  THICKNESS 0.35 ;
  MINENCLOSEDAREA 0.14 ;

  EDGECAPACITANCE 37.759E-6 ;
  CAPACITANCE CPERSQDIST 16.9423E-6 ;
  RESISTANCE RPERSQ 0.125 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met2

# ******** Layer via2, type routing, number 44 **************
LAYER via2
  TYPE CUT ;
  WIDTH 0.2 ;                   # Via2 1
  SPACING 0.2 ;                 # Via2 2
  ENCLOSURE BELOW 0.04 0.085 ;  # Via2 4
  ENCLOSURE ABOVE 0.065 0.065 ; # Met3 4
  RESISTANCE 3.41 ;
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 0.68 ;
  OFFSET 0.34 ;

  WIDTH 0.3 ;              # Met3 1
  # SPACING 0.3 ;          # Met3 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.3
     WIDTH 3 0.4 ;
  AREA 0.24 ;              # Met3 6
  THICKNESS 0.8 ;

  EDGECAPACITANCE 40.989E-6 ;
  CAPACITANCE CPERSQDIST 12.3729E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met3

LAYER via3
  TYPE CUT ;
  WIDTH 0.2 ;                   # Via3 1
  SPACING 0.2 ;                 # Via3 2
  ENCLOSURE BELOW 0.06 0.09 ;   # Via3 4 / Via3 5
  ENCLOSURE ABOVE 0.065 0.065 ; # Met4 3
  RESISTANCE 3.41 ;
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.92 ;
  OFFSET 0.46 ;

  WIDTH 0.3 ;             # Met4 1
  # SPACING  0.3 ;             # Met4 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.3
     WIDTH 3 0.4 ;
  AREA 0.24 ;            # Met4 4a

  THICKNESS 0.8 ;

  EDGECAPACITANCE 36.676E-6 ;
  CAPACITANCE CPERSQDIST 8.41537E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  MAXIMUMDENSITY 70 ;
  DENSITYCHECKWINDOW 700 700 ;
  DENSITYCHECKSTEP 70 ;
END met4

LAYER via4
  TYPE CUT ;

  WIDTH 0.8 ;                 # Via4 1
  SPACING 0.8 ;               # Via4 2
  ENCLOSURE BELOW 0.19 0.19 ; # Via4 4
  ENCLOSURE ABOVE 0.31 0.31 ; # Met5 3
  RESISTANCE 0.38 ;
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 2.49 ; # mA per via Iavg_max at Tj = 90oC
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 3.4 ;
  OFFSET 1.7 ;

  WIDTH 1.6 ;            # Met5 1
  #SPACING  1.6 ;        # Met5 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 1.6 ;
  AREA 4 ;               # Met5 4

  THICKNESS 1.2 ;

  EDGECAPACITANCE 38.851E-6 ;
  CAPACITANCE CPERSQDIST 6.32063E-6 ;
  RESISTANCE RPERSQ 0.0285 ;
  DCCURRENTDENSITY AVERAGE 10.17 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 22.34 ; # mA/um Irms_max at Tj = 90oC

  ANTENNAMODEL OXIDE1 ;
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met5


### Routing via cells section   ###
# Plus via rule, metals are along the prefered direction
VIA L1M1_PR DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIARULE L1M1_PR GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.03 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR

# Plus via rule, metals are along the non prefered direction
VIA L1M1_PR_R DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIARULE L1M1_PR_R GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.03 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA L1M1_PR_M DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIARULE L1M1_PR_M GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.03 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA L1M1_PR_MR DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIARULE L1M1_PR_MR GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.03 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_MR

# Centered via rule, we really do not want to use it
VIA L1M1_PR_C DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIARULE L1M1_PR_C GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_C

# Plus via rule, metals are along the prefered direction
VIA M1M2_PR DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.13 0.16 0.13 ;
  LAYER met2 ;
  RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIARULE M1M2_PR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR

# Plus via rule, metals are along the non prefered direction
VIA M1M2_PR_R DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.13 -0.16 0.13 0.16 ;
  LAYER met2 ;
  RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIARULE M1M2_PR_R GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M1M2_PR_M DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.13 0.16 0.13 ;
  LAYER met2 ;
  RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIARULE M1M2_PR_M GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M1M2_PR_MR DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.13 -0.16 0.13 0.16 ;
  LAYER met2 ;
  RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIARULE M1M2_PR_MR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_MR

# Centered via rule, we really do not want to use it
VIA M1M2_PR_C DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.16 0.16 0.16 ;
  LAYER met2 ;
  RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIARULE M1M2_PR_C GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_C

# Plus via rule, metals are along the prefered direction
VIA M2M3_PR DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.185 0.14 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIARULE M2M3_PR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR

# Plus via rule, metals are along the non prefered direction
VIA M2M3_PR_R DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.14 0.185 0.14 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIARULE M2M3_PR_R GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.04 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M2M3_PR_M DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.185 0.14 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIARULE M2M3_PR_M GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M2M3_PR_MR DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.14 0.185 0.14 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIARULE M2M3_PR_MR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.04 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_MR

# Centered via rule, we really do not want to use it
VIA M2M3_PR_C DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.185 0.185 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIARULE M2M3_PR_C GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_C

# Plus via rule, metals are along the prefered direction
VIA M3M4_PR DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.16 0.19 0.16 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIARULE M3M4_PR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.06 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR

# Plus via rule, metals are along the non prefered direction
VIA M3M4_PR_R DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.16 -0.19 0.16 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIARULE M3M4_PR_R GENERATE
  LAYER met3 ;
  ENCLOSURE 0.06 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M3M4_PR_M DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.16 0.19 0.16 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIARULE M3M4_PR_M GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.06 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M3M4_PR_MR DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.16 -0.19 0.16 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIARULE M3M4_PR_MR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.06 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_MR

# Centered via rule, we really do not want to use it
VIA M3M4_PR_C DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.19 0.19 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIARULE M3M4_PR_C GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_C

# Plus via rule, metals are along the prefered direction
VIA M4M5_PR DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIARULE M4M5_PR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR

# Plus via rule, metals are along the non prefered direction
VIA M4M5_PR_R DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIARULE M4M5_PR_R GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M4M5_PR_M DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIARULE M4M5_PR_M GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M4M5_PR_MR DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIARULE M4M5_PR_MR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_MR

# Centered via rule, we really do not want to use it
VIA M4M5_PR_C DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

VIARULE M4M5_PR_C GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_C
###  end of single via cells   ###

END LIBRARY
VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_hd__a2bb2o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.910 0.995 1.240 1.615 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.410 0.995 1.700 1.375 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 3.280 0.765 3.540 1.655 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.600 1.355 3.080 1.655 ;
        RECT 2.820 0.765 3.080 1.355 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 0.925 1.015 ;
        RECT 0.005 0.105 3.590 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.525 0.345 2.465 ;
        RECT 0.085 0.810 0.260 1.525 ;
        RECT 0.085 0.255 0.345 0.810 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.515 2.235 0.845 2.635 ;
        RECT 1.990 2.370 2.245 2.465 ;
        RECT 1.105 2.200 2.245 2.370 ;
        RECT 2.415 2.255 2.745 2.425 ;
        RECT 1.105 1.975 1.275 2.200 ;
        RECT 0.515 1.805 1.275 1.975 ;
        RECT 1.990 2.065 2.245 2.200 ;
        RECT 0.515 1.325 0.685 1.805 ;
        RECT 1.540 1.715 1.710 1.905 ;
        RECT 1.990 1.895 2.400 2.065 ;
        RECT 1.540 1.545 2.060 1.715 ;
        RECT 0.430 0.995 0.685 1.325 ;
        RECT 1.890 0.825 2.060 1.545 ;
        RECT 1.180 0.655 2.060 0.825 ;
        RECT 2.230 0.870 2.400 1.895 ;
        RECT 2.575 2.005 2.745 2.255 ;
        RECT 2.915 2.175 3.165 2.635 ;
        RECT 3.335 2.005 3.515 2.465 ;
        RECT 2.575 1.835 3.515 2.005 ;
        RECT 2.230 0.700 2.580 0.870 ;
        RECT 0.515 0.085 0.945 0.530 ;
        RECT 1.180 0.255 1.350 0.655 ;
        RECT 1.520 0.085 2.240 0.485 ;
        RECT 2.410 0.255 2.580 0.700 ;
        RECT 3.155 0.085 3.555 0.595 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__a2bb2o_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a2bb2o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.345 0.995 1.675 1.615 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.845 0.995 2.135 1.375 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 3.730 0.765 3.990 1.655 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 3.050 1.355 3.530 1.655 ;
        RECT 3.270 0.765 3.530 1.355 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.785 1.360 1.015 ;
        RECT 0.015 0.105 4.040 0.785 ;
        RECT 0.125 -0.085 0.295 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.525 0.780 2.465 ;
        RECT 0.525 0.810 0.695 1.525 ;
        RECT 0.525 0.255 0.780 0.810 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.185 1.445 0.355 2.635 ;
        RECT 0.950 2.235 1.280 2.635 ;
        RECT 2.500 2.370 2.670 2.465 ;
        RECT 1.540 2.200 2.670 2.370 ;
        RECT 2.875 2.255 3.205 2.425 ;
        RECT 1.540 1.975 1.710 2.200 ;
        RECT 0.950 1.805 1.710 1.975 ;
        RECT 2.440 2.065 2.670 2.200 ;
        RECT 0.950 1.325 1.120 1.805 ;
        RECT 1.975 1.715 2.145 1.905 ;
        RECT 2.440 1.895 2.850 2.065 ;
        RECT 1.975 1.545 2.510 1.715 ;
        RECT 0.865 0.995 1.120 1.325 ;
        RECT 0.185 0.085 0.355 0.930 ;
        RECT 2.340 0.825 2.510 1.545 ;
        RECT 1.615 0.655 2.510 0.825 ;
        RECT 2.680 0.870 2.850 1.895 ;
        RECT 3.035 2.005 3.205 2.255 ;
        RECT 3.375 2.175 3.625 2.635 ;
        RECT 3.795 2.005 3.965 2.465 ;
        RECT 3.035 1.835 3.965 2.005 ;
        RECT 2.680 0.700 3.030 0.870 ;
        RECT 0.950 0.085 1.380 0.530 ;
        RECT 1.615 0.255 1.785 0.655 ;
        RECT 1.955 0.085 2.690 0.485 ;
        RECT 2.860 0.255 3.030 0.700 ;
        RECT 3.605 0.085 4.005 0.595 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__a2bb2o_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a2bb2o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.475 1.445 4.965 1.615 ;
        RECT 3.475 1.325 3.645 1.445 ;
        RECT 3.315 1.075 3.645 1.325 ;
        RECT 4.605 1.075 4.965 1.445 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.815 1.075 4.435 1.275 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.445 1.685 1.615 ;
        RECT 0.085 1.075 0.575 1.445 ;
        RECT 1.515 1.245 1.685 1.445 ;
        RECT 1.515 1.075 1.895 1.245 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.805 1.075 1.345 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.915 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 5.275 1.955 5.525 2.465 ;
        RECT 6.115 1.955 6.365 2.465 ;
        RECT 5.275 1.785 6.365 1.955 ;
        RECT 6.115 1.655 6.365 1.785 ;
        RECT 6.115 1.415 6.920 1.655 ;
        RECT 6.610 0.905 6.920 1.415 ;
        RECT 5.235 0.725 6.920 0.905 ;
        RECT 5.235 0.275 5.565 0.725 ;
        RECT 6.075 0.275 6.405 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.135 1.955 0.385 2.465 ;
        RECT 0.555 2.125 0.805 2.635 ;
        RECT 0.975 1.955 1.225 2.465 ;
        RECT 1.395 2.125 1.645 2.635 ;
        RECT 1.815 2.295 2.905 2.465 ;
        RECT 1.815 1.955 2.065 2.295 ;
        RECT 2.655 2.135 2.905 2.295 ;
        RECT 3.175 2.135 3.425 2.635 ;
        RECT 3.595 2.295 4.685 2.465 ;
        RECT 3.595 2.135 3.845 2.295 ;
        RECT 0.135 1.785 2.065 1.955 ;
        RECT 1.855 1.455 2.065 1.785 ;
        RECT 2.235 1.965 2.485 2.125 ;
        RECT 4.015 1.965 4.265 2.125 ;
        RECT 2.235 1.415 2.620 1.965 ;
        RECT 3.135 1.785 4.265 1.965 ;
        RECT 4.435 1.785 4.685 2.295 ;
        RECT 4.855 1.795 5.105 2.635 ;
        RECT 5.695 2.165 5.945 2.635 ;
        RECT 6.535 1.825 6.785 2.635 ;
        RECT 3.135 1.665 3.305 1.785 ;
        RECT 2.955 1.495 3.305 1.665 ;
        RECT 2.235 0.905 2.445 1.415 ;
        RECT 2.955 1.245 3.145 1.495 ;
        RECT 2.615 1.075 3.145 1.245 ;
        RECT 5.135 1.245 5.460 1.615 ;
        RECT 5.135 1.075 6.440 1.245 ;
        RECT 2.955 0.905 3.145 1.075 ;
        RECT 0.175 0.085 0.345 0.895 ;
        RECT 0.515 0.475 0.765 0.905 ;
        RECT 0.935 0.735 2.525 0.905 ;
        RECT 0.935 0.645 1.270 0.735 ;
        RECT 0.515 0.255 1.685 0.475 ;
        RECT 1.855 0.085 2.025 0.555 ;
        RECT 2.195 0.255 2.525 0.735 ;
        RECT 2.955 0.725 4.725 0.905 ;
        RECT 2.695 0.085 3.385 0.555 ;
        RECT 3.555 0.255 3.885 0.725 ;
        RECT 4.055 0.085 4.225 0.555 ;
        RECT 4.395 0.255 4.725 0.725 ;
        RECT 4.895 0.085 5.065 0.895 ;
        RECT 5.735 0.085 5.905 0.555 ;
        RECT 6.575 0.085 6.745 0.555 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 2.450 1.445 2.620 1.615 ;
        RECT 5.230 1.445 5.400 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
      LAYER met1 ;
        RECT 2.390 1.600 2.680 1.645 ;
        RECT 5.170 1.600 5.460 1.645 ;
        RECT 2.390 1.460 5.460 1.600 ;
        RECT 2.390 1.415 2.680 1.460 ;
        RECT 5.170 1.415 5.460 1.460 ;
  END
END sky130_fd_sc_hd__a2bb2o_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a2bb2oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.150 0.995 0.520 1.615 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.725 1.010 1.240 1.275 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.780 0.995 3.070 1.615 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.245 0.995 2.610 1.615 ;
        RECT 2.440 0.425 2.610 0.995 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.215 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.515500 ;
    PORT
      LAYER li1 ;
        RECT 1.420 1.955 1.785 2.465 ;
        RECT 1.420 1.785 1.945 1.955 ;
        RECT 1.775 0.825 1.945 1.785 ;
        RECT 1.775 0.255 2.205 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.095 1.805 0.425 2.635 ;
        RECT 0.875 1.615 1.205 2.465 ;
        RECT 1.955 2.235 2.285 2.465 ;
        RECT 2.115 1.955 2.285 2.235 ;
        RECT 2.455 2.135 2.705 2.635 ;
        RECT 2.875 1.955 3.130 2.465 ;
        RECT 2.115 1.785 3.130 1.955 ;
        RECT 0.875 1.445 1.580 1.615 ;
        RECT 1.410 0.830 1.580 1.445 ;
        RECT 0.095 0.085 0.425 0.825 ;
        RECT 0.595 0.660 1.580 0.830 ;
        RECT 0.595 0.255 0.765 0.660 ;
        RECT 0.935 0.085 1.605 0.490 ;
        RECT 2.795 0.085 3.125 0.825 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__a2bb2oi_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a2bb2oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.310 1.075 4.205 1.275 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.455 1.075 5.435 1.275 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.445 2.030 1.615 ;
        RECT 0.085 1.075 0.710 1.445 ;
        RECT 1.700 1.075 2.030 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.940 1.075 1.480 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140 0.105 5.390 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.621000 ;
    PORT
      LAYER li1 ;
        RECT 2.370 1.660 2.620 2.125 ;
        RECT 2.370 0.905 2.660 1.660 ;
        RECT 1.070 0.725 2.660 0.905 ;
        RECT 1.070 0.645 1.400 0.725 ;
        RECT 2.330 0.255 2.660 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.270 1.955 0.520 2.465 ;
        RECT 0.690 2.135 0.940 2.635 ;
        RECT 1.110 1.955 1.360 2.465 ;
        RECT 1.530 2.135 1.780 2.635 ;
        RECT 1.950 2.295 3.040 2.465 ;
        RECT 1.950 1.955 2.200 2.295 ;
        RECT 0.270 1.785 2.200 1.955 ;
        RECT 2.790 1.795 3.040 2.295 ;
        RECT 3.310 1.965 3.560 2.465 ;
        RECT 3.730 2.135 3.980 2.635 ;
        RECT 4.150 2.295 5.240 2.465 ;
        RECT 4.150 1.965 4.400 2.295 ;
        RECT 3.310 1.785 4.400 1.965 ;
        RECT 4.570 1.615 4.820 2.125 ;
        RECT 2.950 1.445 4.820 1.615 ;
        RECT 4.990 1.455 5.240 2.295 ;
        RECT 2.950 1.325 3.120 1.445 ;
        RECT 2.830 0.995 3.120 1.325 ;
        RECT 2.950 0.905 3.120 0.995 ;
        RECT 0.310 0.085 0.480 0.895 ;
        RECT 0.650 0.475 0.900 0.895 ;
        RECT 2.950 0.725 4.860 0.905 ;
        RECT 0.650 0.255 1.820 0.475 ;
        RECT 1.990 0.085 2.160 0.555 ;
        RECT 2.830 0.085 3.520 0.555 ;
        RECT 3.690 0.255 4.020 0.725 ;
        RECT 4.190 0.085 4.360 0.555 ;
        RECT 4.530 0.255 4.860 0.725 ;
        RECT 5.030 0.085 5.200 0.905 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__a2bb2oi_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a2bb2oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2bb2oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 5.945 1.075 7.320 1.275 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 7.595 1.075 9.045 1.275 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.385 1.445 3.575 1.615 ;
        RECT 1.385 1.285 1.555 1.445 ;
        RECT 0.100 1.075 1.555 1.285 ;
        RECT 3.245 1.075 3.575 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.725 1.075 3.075 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.435 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER li1 ;
        RECT 3.915 1.615 4.165 2.125 ;
        RECT 4.745 1.615 4.965 2.125 ;
        RECT 3.745 1.415 4.965 1.615 ;
        RECT 3.745 0.905 3.915 1.415 ;
        RECT 1.775 0.725 5.045 0.905 ;
        RECT 1.775 0.645 2.995 0.725 ;
        RECT 3.875 0.275 4.205 0.725 ;
        RECT 4.715 0.275 5.045 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.085 1.625 0.425 2.465 ;
        RECT 0.595 1.795 0.805 2.635 ;
        RECT 0.975 1.965 1.215 2.465 ;
        RECT 1.395 2.135 1.645 2.635 ;
        RECT 1.815 1.965 2.065 2.465 ;
        RECT 2.235 2.135 2.485 2.635 ;
        RECT 2.655 1.965 2.905 2.465 ;
        RECT 3.075 2.135 3.325 2.635 ;
        RECT 3.495 2.295 5.465 2.465 ;
        RECT 3.495 1.965 3.745 2.295 ;
        RECT 0.975 1.795 3.745 1.965 ;
        RECT 4.335 1.795 4.575 2.295 ;
        RECT 0.975 1.625 1.215 1.795 ;
        RECT 0.085 1.455 1.215 1.625 ;
        RECT 5.135 1.455 5.465 2.295 ;
        RECT 5.655 1.625 5.985 2.465 ;
        RECT 6.155 1.795 6.365 2.635 ;
        RECT 6.540 1.625 6.780 2.465 ;
        RECT 6.955 1.795 7.205 2.635 ;
        RECT 7.375 2.295 9.310 2.465 ;
        RECT 7.375 1.625 7.625 2.295 ;
        RECT 5.655 1.455 7.625 1.625 ;
        RECT 7.795 1.625 8.045 2.125 ;
        RECT 8.215 1.795 8.465 2.295 ;
        RECT 8.635 1.625 8.885 2.125 ;
        RECT 9.060 1.795 9.310 2.295 ;
        RECT 7.795 1.455 9.575 1.625 ;
        RECT 4.085 1.075 5.725 1.245 ;
        RECT 5.555 0.905 5.725 1.075 ;
        RECT 9.215 0.905 9.575 1.455 ;
        RECT 0.175 0.085 0.345 0.895 ;
        RECT 0.515 0.725 1.605 0.905 ;
        RECT 5.555 0.735 9.575 0.905 ;
        RECT 0.515 0.255 0.845 0.725 ;
        RECT 1.015 0.085 1.185 0.555 ;
        RECT 1.355 0.475 1.605 0.725 ;
        RECT 6.075 0.725 8.925 0.735 ;
        RECT 1.355 0.255 3.365 0.475 ;
        RECT 3.535 0.085 3.705 0.555 ;
        RECT 4.375 0.085 4.545 0.555 ;
        RECT 5.215 0.085 5.905 0.555 ;
        RECT 6.075 0.255 6.405 0.725 ;
        RECT 6.575 0.085 6.745 0.555 ;
        RECT 6.915 0.255 7.245 0.725 ;
        RECT 7.415 0.085 7.585 0.555 ;
        RECT 7.755 0.255 8.085 0.725 ;
        RECT 8.255 0.085 8.425 0.555 ;
        RECT 8.595 0.255 8.925 0.725 ;
        RECT 9.095 0.085 9.265 0.555 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
  END
END sky130_fd_sc_hd__a2bb2oi_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a21bo_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21bo_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.750 0.995 2.175 1.615 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.370 0.995 2.630 1.615 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.325 0.335 1.665 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 3.300 0.265 3.580 2.455 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 0.850 0.785 3.675 1.015 ;
        RECT 0.345 0.105 3.675 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.105 2.045 0.345 2.435 ;
        RECT 0.515 2.225 0.865 2.635 ;
        RECT 0.105 1.845 0.855 2.045 ;
        RECT 0.515 1.165 0.855 1.845 ;
        RECT 1.035 1.345 1.365 2.455 ;
        RECT 1.535 1.985 1.715 2.455 ;
        RECT 1.885 2.155 2.215 2.635 ;
        RECT 2.390 1.985 2.560 2.455 ;
        RECT 1.535 1.785 2.560 1.985 ;
        RECT 2.825 1.495 3.110 2.635 ;
        RECT 0.515 0.265 0.745 1.165 ;
        RECT 1.035 1.045 1.580 1.345 ;
        RECT 0.945 0.085 1.190 0.865 ;
        RECT 1.360 0.815 1.580 1.045 ;
        RECT 2.840 0.815 3.100 1.325 ;
        RECT 1.360 0.625 3.100 0.815 ;
        RECT 1.360 0.265 1.790 0.625 ;
        RECT 2.370 0.085 3.100 0.455 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__a21bo_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a21bo_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21bo_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.685 0.995 3.100 1.615 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.270 0.995 3.560 1.615 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.070 1.035 1.525 1.325 ;
        RECT 1.330 0.995 1.525 1.035 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.655 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER li1 ;
        RECT 0.595 2.005 0.850 2.425 ;
        RECT 0.150 1.835 0.850 2.005 ;
        RECT 0.150 0.885 0.380 1.835 ;
        RECT 0.150 0.715 0.850 0.885 ;
        RECT 0.520 0.315 0.850 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.090 2.255 0.425 2.635 ;
        RECT 1.040 2.275 1.370 2.635 ;
        RECT 1.975 2.105 2.225 2.465 ;
        RECT 1.115 1.895 2.225 2.105 ;
        RECT 1.115 1.665 1.285 1.895 ;
        RECT 0.570 1.495 1.285 1.665 ;
        RECT 1.455 1.555 1.865 1.725 ;
        RECT 0.570 1.075 0.900 1.495 ;
        RECT 1.695 1.325 1.865 1.555 ;
        RECT 2.055 1.675 2.225 1.895 ;
        RECT 2.395 2.015 2.725 2.465 ;
        RECT 2.895 2.185 3.065 2.635 ;
        RECT 3.235 2.015 3.565 2.465 ;
        RECT 2.395 1.845 3.565 2.015 ;
        RECT 2.055 1.505 2.515 1.675 ;
        RECT 1.695 0.995 2.175 1.325 ;
        RECT 0.090 0.085 0.345 0.545 ;
        RECT 1.020 0.085 1.220 0.865 ;
        RECT 1.695 0.825 1.865 0.995 ;
        RECT 1.455 0.655 1.865 0.825 ;
        RECT 2.345 0.825 2.515 1.505 ;
        RECT 2.345 0.635 2.740 0.825 ;
        RECT 1.975 0.085 2.305 0.465 ;
        RECT 3.235 0.085 3.565 0.825 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__a21bo_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a21bo_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21bo_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.590 1.010 4.955 1.360 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.245 1.595 5.390 1.765 ;
        RECT 4.245 1.275 4.420 1.595 ;
        RECT 4.025 1.010 4.420 1.275 ;
        RECT 5.220 1.290 5.390 1.595 ;
        RECT 5.220 1.055 5.700 1.290 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.500 1.010 0.830 1.625 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.080 0.105 5.915 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER li1 ;
        RECT 1.000 1.595 2.410 1.765 ;
        RECT 1.000 0.785 1.235 1.595 ;
        RECT 1.000 0.615 2.340 0.785 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.105 2.105 0.550 2.465 ;
        RECT 0.720 2.275 1.050 2.635 ;
        RECT 1.580 2.275 1.910 2.635 ;
        RECT 2.435 2.275 2.770 2.635 ;
        RECT 3.055 2.210 4.065 2.380 ;
        RECT 4.235 2.275 4.565 2.635 ;
        RECT 5.075 2.275 5.405 2.635 ;
        RECT 0.105 1.935 2.870 2.105 ;
        RECT 0.105 1.795 0.565 1.935 ;
        RECT 0.105 0.840 0.330 1.795 ;
        RECT 2.700 1.525 2.870 1.935 ;
        RECT 3.055 1.695 3.225 2.210 ;
        RECT 3.885 2.105 4.065 2.210 ;
        RECT 3.885 1.935 5.825 2.105 ;
        RECT 2.700 1.355 3.305 1.525 ;
        RECT 1.405 1.185 2.530 1.325 ;
        RECT 1.405 0.995 2.810 1.185 ;
        RECT 2.995 0.995 3.305 1.355 ;
        RECT 0.105 0.255 0.540 0.840 ;
        RECT 2.640 0.800 2.810 0.995 ;
        RECT 3.475 0.840 3.645 1.805 ;
        RECT 3.885 1.445 4.065 1.935 ;
        RECT 5.570 1.460 5.825 1.935 ;
        RECT 2.640 0.785 3.010 0.800 ;
        RECT 3.475 0.785 4.965 0.840 ;
        RECT 2.640 0.670 4.965 0.785 ;
        RECT 2.640 0.615 3.645 0.670 ;
        RECT 0.710 0.085 1.050 0.445 ;
        RECT 1.580 0.085 1.910 0.445 ;
        RECT 2.515 0.085 3.285 0.445 ;
        RECT 3.475 0.255 3.645 0.615 ;
        RECT 3.855 0.085 4.185 0.445 ;
        RECT 4.685 0.405 4.965 0.670 ;
        RECT 5.545 0.085 5.825 0.885 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
END sky130_fd_sc_hd__a21bo_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a21boi_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.780 0.765 2.170 1.615 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.340 0.765 2.615 1.435 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.470 1.200 0.895 1.955 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.755 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.392200 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.655 1.305 2.465 ;
        RECT 1.065 1.200 1.610 1.655 ;
        RECT 1.315 0.255 1.610 1.200 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.095 2.085 0.355 2.465 ;
        RECT 0.525 2.175 0.855 2.635 ;
        RECT 0.095 1.030 0.300 2.085 ;
        RECT 1.475 2.005 1.805 2.465 ;
        RECT 1.975 2.175 2.165 2.635 ;
        RECT 2.335 2.005 2.665 2.465 ;
        RECT 1.475 1.825 2.665 2.005 ;
        RECT 0.095 0.780 1.145 1.030 ;
        RECT 0.095 0.280 0.380 0.780 ;
        RECT 0.550 0.085 1.145 0.610 ;
        RECT 2.335 0.085 2.665 0.595 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__a21boi_0

#--------EOF---------

MACRO sky130_fd_sc_hd__a21boi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.760 0.995 2.155 1.345 ;
        RECT 1.945 0.375 2.155 0.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.350 0.995 2.640 1.345 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.975 0.335 1.665 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.785 0.785 2.745 1.015 ;
        RECT 0.295 0.105 2.745 0.785 ;
        RECT 0.295 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.551000 ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.345 1.375 2.455 ;
        RECT 1.045 1.045 1.580 1.345 ;
        RECT 1.335 0.795 1.580 1.045 ;
        RECT 1.335 0.265 1.765 0.795 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.095 2.045 0.355 2.435 ;
        RECT 0.525 2.225 0.855 2.635 ;
        RECT 0.095 1.845 0.855 2.045 ;
        RECT 0.515 1.165 0.855 1.845 ;
        RECT 1.545 1.725 1.735 2.455 ;
        RECT 1.905 1.905 2.235 2.635 ;
        RECT 2.415 1.725 2.585 2.455 ;
        RECT 1.545 1.525 2.585 1.725 ;
        RECT 0.515 0.715 0.745 1.165 ;
        RECT 0.365 0.265 0.745 0.715 ;
        RECT 0.925 0.085 1.155 0.865 ;
        RECT 2.325 0.085 2.655 0.815 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__a21boi_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a21boi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.605 0.995 3.215 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.100 1.495 3.675 1.675 ;
        RECT 2.100 1.245 2.425 1.495 ;
        RECT 2.095 1.075 2.425 1.245 ;
        RECT 3.385 1.295 3.675 1.495 ;
        RECT 3.385 1.035 3.795 1.295 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.120 0.765 0.425 1.805 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.700 0.785 4.030 1.015 ;
        RECT 0.175 0.105 4.030 0.785 ;
        RECT 0.175 0.085 0.320 0.105 ;
        RECT 0.150 -0.085 0.320 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.627500 ;
    PORT
      LAYER li1 ;
        RECT 1.520 0.785 1.715 2.115 ;
        RECT 1.520 0.615 3.060 0.785 ;
        RECT 1.520 0.255 1.720 0.615 ;
        RECT 2.730 0.255 3.060 0.615 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.095 2.080 0.425 2.635 ;
        RECT 1.045 2.285 2.215 2.465 ;
        RECT 0.595 1.285 0.855 2.265 ;
        RECT 1.045 1.795 1.350 2.285 ;
        RECT 1.885 2.025 2.215 2.285 ;
        RECT 2.385 2.195 2.555 2.635 ;
        RECT 2.810 2.105 2.980 2.465 ;
        RECT 3.160 2.275 3.490 2.635 ;
        RECT 3.660 2.105 3.920 2.465 ;
        RECT 2.810 2.025 3.920 2.105 ;
        RECT 1.885 1.855 3.920 2.025 ;
        RECT 0.595 1.070 1.325 1.285 ;
        RECT 0.595 0.530 0.795 1.070 ;
        RECT 0.265 0.360 0.795 0.530 ;
        RECT 0.985 0.085 1.225 0.885 ;
        RECT 1.940 0.085 2.270 0.445 ;
        RECT 3.635 0.085 3.930 0.865 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__a21boi_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a21boi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21boi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.545 1.065 4.970 1.310 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.030 1.480 6.450 1.705 ;
        RECT 3.030 1.065 3.375 1.480 ;
        RECT 5.205 1.075 6.450 1.480 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.145 1.075 0.650 1.615 ;
        RECT 0.480 0.995 0.650 1.075 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.695 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.288000 ;
    PORT
      LAYER li1 ;
        RECT 1.560 1.705 2.725 2.035 ;
        RECT 1.560 1.585 2.860 1.705 ;
        RECT 2.570 0.895 2.860 1.585 ;
        RECT 2.570 0.865 4.885 0.895 ;
        RECT 1.275 0.695 4.885 0.865 ;
        RECT 1.275 0.615 2.325 0.695 ;
        RECT 3.255 0.675 4.885 0.695 ;
        RECT 1.275 0.370 1.465 0.615 ;
        RECT 2.135 0.255 2.325 0.615 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.125 2.005 0.455 2.465 ;
        RECT 0.625 2.175 0.885 2.635 ;
        RECT 1.160 2.215 3.095 2.465 ;
        RECT 3.265 2.275 3.595 2.635 ;
        RECT 4.125 2.275 4.455 2.635 ;
        RECT 0.125 1.785 0.990 2.005 ;
        RECT 1.160 1.795 1.355 2.215 ;
        RECT 1.935 2.205 3.095 2.215 ;
        RECT 2.895 2.105 3.095 2.205 ;
        RECT 4.625 2.105 4.815 2.465 ;
        RECT 4.985 2.275 5.315 2.635 ;
        RECT 5.485 2.105 5.665 2.465 ;
        RECT 5.845 2.275 6.175 2.635 ;
        RECT 6.345 2.105 6.605 2.465 ;
        RECT 2.895 1.875 6.605 2.105 ;
        RECT 0.820 1.345 0.990 1.785 ;
        RECT 0.820 1.035 2.400 1.345 ;
        RECT 0.820 0.795 1.105 1.035 ;
        RECT 0.090 0.615 1.105 0.795 ;
        RECT 5.055 0.735 6.175 0.905 ;
        RECT 0.090 0.255 0.445 0.615 ;
        RECT 0.720 0.085 1.105 0.445 ;
        RECT 1.635 0.085 1.965 0.445 ;
        RECT 2.495 0.085 3.085 0.525 ;
        RECT 5.055 0.505 5.315 0.735 ;
        RECT 3.265 0.255 5.315 0.505 ;
        RECT 5.485 0.085 5.675 0.565 ;
        RECT 5.845 0.255 6.175 0.735 ;
        RECT 6.345 0.085 6.605 0.885 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
  END
END sky130_fd_sc_hd__a21boi_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a21o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.660 1.015 2.185 1.325 ;
        RECT 1.955 0.375 2.185 1.015 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.365 0.995 2.665 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.015 1.480 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.105 2.745 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.265 0.355 2.455 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.525 1.905 0.865 2.635 ;
        RECT 1.045 1.725 1.315 2.455 ;
        RECT 0.545 1.505 1.315 1.725 ;
        RECT 1.495 1.745 1.725 2.455 ;
        RECT 1.895 1.925 2.225 2.635 ;
        RECT 2.395 1.745 2.655 2.455 ;
        RECT 1.495 1.505 2.655 1.745 ;
        RECT 0.545 0.835 0.835 1.505 ;
        RECT 0.545 0.635 1.775 0.835 ;
        RECT 0.615 0.085 1.285 0.455 ;
        RECT 1.465 0.265 1.775 0.635 ;
        RECT 2.365 0.085 2.655 0.815 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__a21o_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a21o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.240 0.365 2.620 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.810 0.750 3.125 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.465 0.995 1.790 1.410 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.175 0.105 3.215 1.015 ;
        RECT 0.175 0.085 0.320 0.105 ;
        RECT 0.150 -0.085 0.320 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER li1 ;
        RECT 0.555 0.825 0.785 2.465 ;
        RECT 0.555 0.635 0.955 0.825 ;
        RECT 0.765 0.255 0.955 0.635 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.095 1.665 0.385 2.635 ;
        RECT 0.955 2.220 1.285 2.635 ;
        RECT 1.475 1.920 1.790 2.465 ;
        RECT 0.955 1.690 1.790 1.920 ;
        RECT 1.960 1.935 2.185 2.465 ;
        RECT 2.355 2.125 2.685 2.635 ;
        RECT 2.855 1.935 3.075 2.465 ;
        RECT 0.955 0.995 1.295 1.690 ;
        RECT 1.960 1.670 3.075 1.935 ;
        RECT 1.125 0.825 1.295 0.995 ;
        RECT 1.125 0.655 1.865 0.825 ;
        RECT 0.265 0.085 0.595 0.465 ;
        RECT 1.125 0.085 1.455 0.445 ;
        RECT 1.675 0.255 1.865 0.655 ;
        RECT 2.805 0.085 3.135 0.565 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__a21o_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a21o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.990 1.010 4.515 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.645 1.510 4.935 1.680 ;
        RECT 3.645 1.275 3.820 1.510 ;
        RECT 3.425 1.010 3.820 1.275 ;
        RECT 4.685 1.290 4.935 1.510 ;
        RECT 4.685 1.055 5.100 1.290 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.395 0.995 2.705 1.525 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.315 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER li1 ;
        RECT 0.625 1.755 0.795 2.185 ;
        RECT 1.485 1.755 1.735 2.185 ;
        RECT 0.145 1.585 1.735 1.755 ;
        RECT 0.145 0.785 0.630 1.585 ;
        RECT 0.145 0.615 1.735 0.785 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.115 1.935 0.445 2.635 ;
        RECT 0.975 1.935 1.305 2.635 ;
        RECT 1.915 1.515 2.165 2.635 ;
        RECT 2.455 2.295 3.465 2.465 ;
        RECT 2.455 1.695 2.625 2.295 ;
        RECT 0.800 0.995 2.205 1.325 ;
        RECT 2.035 0.785 2.205 0.995 ;
        RECT 2.875 0.840 3.045 2.125 ;
        RECT 3.285 2.020 3.465 2.295 ;
        RECT 3.635 2.275 3.965 2.635 ;
        RECT 4.135 2.020 4.305 2.465 ;
        RECT 4.475 2.275 4.805 2.635 ;
        RECT 5.030 2.020 5.360 2.395 ;
        RECT 3.285 1.850 5.360 2.020 ;
        RECT 3.285 1.445 3.465 1.850 ;
        RECT 5.105 1.460 5.360 1.850 ;
        RECT 2.875 0.785 4.365 0.840 ;
        RECT 2.035 0.670 4.365 0.785 ;
        RECT 2.035 0.615 3.045 0.670 ;
        RECT 0.105 0.085 0.445 0.445 ;
        RECT 0.975 0.085 1.305 0.445 ;
        RECT 1.910 0.085 2.685 0.445 ;
        RECT 2.875 0.255 3.045 0.615 ;
        RECT 3.255 0.085 3.585 0.445 ;
        RECT 4.085 0.405 4.365 0.670 ;
        RECT 4.945 0.085 5.225 0.885 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__a21o_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a21oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.850 0.995 1.265 1.325 ;
        RECT 1.035 0.375 1.265 0.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.445 0.995 1.740 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.675 0.335 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.105 1.835 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.447000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.685 0.370 2.455 ;
        RECT 0.095 1.495 0.680 1.685 ;
        RECT 0.505 0.825 0.680 1.495 ;
        RECT 0.505 0.645 0.835 0.825 ;
        RECT 0.610 0.265 0.835 0.645 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.540 2.025 0.870 2.455 ;
        RECT 1.040 2.195 1.235 2.635 ;
        RECT 1.415 2.025 1.745 2.455 ;
        RECT 0.540 1.855 1.745 2.025 ;
        RECT 0.850 1.525 1.745 1.855 ;
        RECT 0.110 0.085 0.440 0.475 ;
        RECT 1.445 0.085 1.745 0.815 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__a21oi_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a21oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.815 0.995 1.425 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 1.495 1.930 1.675 ;
        RECT 0.145 1.035 0.645 1.495 ;
        RECT 1.605 1.245 1.930 1.495 ;
        RECT 1.605 1.075 1.935 1.245 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.800 0.995 3.075 1.625 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.215 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.627500 ;
    PORT
      LAYER li1 ;
        RECT 2.315 0.785 2.615 2.115 ;
        RECT 0.955 0.615 2.615 0.785 ;
        RECT 0.955 0.255 1.300 0.615 ;
        RECT 2.295 0.255 2.615 0.615 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.110 2.105 0.370 2.465 ;
        RECT 0.540 2.275 0.870 2.635 ;
        RECT 1.050 2.105 1.220 2.465 ;
        RECT 1.475 2.195 1.645 2.635 ;
        RECT 1.815 2.285 3.090 2.465 ;
        RECT 0.110 2.025 1.220 2.105 ;
        RECT 1.815 2.025 2.145 2.285 ;
        RECT 0.110 1.855 2.145 2.025 ;
        RECT 2.785 1.795 3.090 2.285 ;
        RECT 0.100 0.085 0.395 0.865 ;
        RECT 1.760 0.085 2.090 0.445 ;
        RECT 2.795 0.085 3.125 0.825 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__a21oi_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a21oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a21oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 2.565 1.065 4.000 1.310 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 2.050 1.480 5.470 1.705 ;
        RECT 2.050 1.065 2.395 1.480 ;
        RECT 4.225 1.075 5.470 1.480 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.035 1.430 1.415 ;
        RECT 0.090 0.995 0.400 1.035 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.715 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.288000 ;
    PORT
      LAYER li1 ;
        RECT 0.580 1.705 1.745 2.035 ;
        RECT 0.580 1.585 1.880 1.705 ;
        RECT 1.600 0.895 1.880 1.585 ;
        RECT 1.600 0.865 3.905 0.895 ;
        RECT 0.595 0.695 3.905 0.865 ;
        RECT 0.595 0.615 1.645 0.695 ;
        RECT 2.275 0.675 3.905 0.695 ;
        RECT 0.595 0.370 0.785 0.615 ;
        RECT 1.455 0.255 1.645 0.615 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.180 2.215 2.115 2.465 ;
        RECT 2.285 2.275 2.615 2.635 ;
        RECT 0.180 1.795 0.375 2.215 ;
        RECT 0.955 2.205 2.115 2.215 ;
        RECT 1.915 2.105 2.115 2.205 ;
        RECT 2.785 2.105 2.975 2.465 ;
        RECT 3.145 2.275 3.475 2.635 ;
        RECT 3.645 2.105 3.835 2.465 ;
        RECT 4.005 2.275 4.335 2.635 ;
        RECT 4.505 2.105 4.685 2.465 ;
        RECT 4.865 2.275 5.195 2.635 ;
        RECT 5.365 2.105 5.625 2.465 ;
        RECT 1.915 1.875 5.625 2.105 ;
        RECT 0.090 0.085 0.425 0.805 ;
        RECT 4.075 0.735 5.195 0.905 ;
        RECT 0.955 0.085 1.285 0.445 ;
        RECT 1.835 0.085 2.115 0.525 ;
        RECT 4.075 0.505 4.335 0.735 ;
        RECT 2.285 0.255 4.335 0.505 ;
        RECT 4.505 0.085 4.695 0.565 ;
        RECT 4.865 0.255 5.195 0.735 ;
        RECT 5.365 0.085 5.625 0.885 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
END sky130_fd_sc_hd__a21oi_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a22o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.075 1.815 1.285 ;
        RECT 1.485 0.675 1.695 1.075 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.040 2.395 1.345 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.765 1.075 1.240 1.285 ;
        RECT 1.020 0.675 1.240 1.075 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.575 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.215 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 2.875 1.785 3.135 2.465 ;
        RECT 2.965 0.585 3.135 1.785 ;
        RECT 2.875 0.255 3.135 0.585 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.090 2.245 0.425 2.465 ;
        RECT 1.430 2.255 1.785 2.635 ;
        RECT 0.090 1.625 0.345 2.245 ;
        RECT 0.595 2.085 0.825 2.125 ;
        RECT 1.955 2.085 2.205 2.465 ;
        RECT 0.595 1.885 2.205 2.085 ;
        RECT 0.595 1.795 0.780 1.885 ;
        RECT 1.370 1.875 2.205 1.885 ;
        RECT 2.455 1.855 2.705 2.635 ;
        RECT 0.935 1.685 1.265 1.715 ;
        RECT 0.935 1.625 2.735 1.685 ;
        RECT 0.090 1.515 2.795 1.625 ;
        RECT 0.090 1.455 1.265 1.515 ;
        RECT 2.595 1.480 2.795 1.515 ;
        RECT 2.625 0.905 2.795 1.480 ;
        RECT 0.090 0.085 0.545 0.850 ;
        RECT 2.525 0.785 2.795 0.905 ;
        RECT 1.950 0.740 2.795 0.785 ;
        RECT 1.950 0.615 2.705 0.740 ;
        RECT 1.950 0.465 2.120 0.615 ;
        RECT 0.820 0.255 2.120 0.465 ;
        RECT 2.375 0.085 2.705 0.445 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__a22o_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a22o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.510 1.075 1.840 1.285 ;
        RECT 1.510 0.675 1.720 1.075 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.010 1.075 2.415 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.765 1.075 1.240 1.285 ;
        RECT 1.020 0.675 1.240 1.075 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.575 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.670 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 2.900 1.785 3.160 2.465 ;
        RECT 2.990 0.585 3.160 1.785 ;
        RECT 2.900 0.255 3.160 0.585 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.095 2.295 1.265 2.465 ;
        RECT 0.095 1.625 0.425 2.295 ;
        RECT 0.935 2.255 1.265 2.295 ;
        RECT 1.455 2.215 1.810 2.635 ;
        RECT 0.595 2.035 0.825 2.125 ;
        RECT 1.980 2.035 2.230 2.465 ;
        RECT 0.595 1.795 2.230 2.035 ;
        RECT 2.400 1.875 2.730 2.635 ;
        RECT 0.095 1.455 2.815 1.625 ;
        RECT 2.645 0.905 2.815 1.455 ;
        RECT 3.330 1.445 3.500 2.635 ;
        RECT 0.095 0.085 0.545 0.850 ;
        RECT 1.975 0.735 2.815 0.905 ;
        RECT 1.975 0.505 2.145 0.735 ;
        RECT 0.820 0.255 2.145 0.505 ;
        RECT 2.355 0.085 2.685 0.565 ;
        RECT 3.330 0.085 3.500 0.985 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__a22o_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a22o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.900 1.075 5.395 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.350 1.445 5.735 1.615 ;
        RECT 4.350 1.075 4.680 1.445 ;
        RECT 5.565 1.275 5.735 1.445 ;
        RECT 5.565 1.075 6.355 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.125 1.075 3.680 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.420 1.445 4.180 1.615 ;
        RECT 2.420 1.075 2.955 1.445 ;
        RECT 3.850 1.075 4.180 1.445 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.070 0.105 6.240 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.640 1.615 0.890 2.465 ;
        RECT 1.480 1.615 1.730 2.465 ;
        RECT 0.085 1.445 1.730 1.615 ;
        RECT 0.085 0.905 0.370 1.445 ;
        RECT 0.085 0.725 1.770 0.905 ;
        RECT 0.600 0.265 0.930 0.725 ;
        RECT 1.440 0.255 1.770 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.220 1.825 0.470 2.635 ;
        RECT 1.060 1.795 1.310 2.635 ;
        RECT 1.900 2.125 2.150 2.635 ;
        RECT 2.420 2.295 4.430 2.465 ;
        RECT 2.420 2.125 2.670 2.295 ;
        RECT 3.260 2.125 3.510 2.295 ;
        RECT 2.840 1.955 3.090 2.125 ;
        RECT 3.680 1.955 3.930 2.125 ;
        RECT 1.900 1.785 3.930 1.955 ;
        RECT 4.100 1.955 4.430 2.295 ;
        RECT 4.600 2.125 4.850 2.635 ;
        RECT 5.020 1.955 5.270 2.465 ;
        RECT 5.440 2.125 5.690 2.635 ;
        RECT 5.905 1.955 6.110 2.465 ;
        RECT 4.100 1.785 6.110 1.955 ;
        RECT 1.900 1.275 2.230 1.785 ;
        RECT 5.905 1.455 6.110 1.785 ;
        RECT 0.540 1.075 2.230 1.275 ;
        RECT 1.940 0.905 2.230 1.075 ;
        RECT 1.940 0.735 5.310 0.905 ;
        RECT 3.170 0.645 3.605 0.735 ;
        RECT 4.935 0.645 5.310 0.735 ;
        RECT 0.260 0.085 0.430 0.555 ;
        RECT 1.100 0.085 1.270 0.555 ;
        RECT 1.940 0.085 2.630 0.555 ;
        RECT 2.800 0.255 3.970 0.475 ;
        RECT 4.185 0.085 4.355 0.555 ;
        RECT 5.480 0.475 5.730 0.895 ;
        RECT 4.560 0.255 5.730 0.475 ;
        RECT 5.900 0.085 6.070 0.895 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
END sky130_fd_sc_hd__a22o_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a22oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.490 1.075 1.840 1.275 ;
        RECT 1.490 0.675 1.700 1.075 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.010 0.995 2.335 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.765 1.075 1.240 1.275 ;
        RECT 0.990 0.675 1.240 1.075 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.765 0.575 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.755 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.858000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 2.295 1.265 2.465 ;
        RECT 0.095 1.625 0.425 2.295 ;
        RECT 0.935 2.255 1.265 2.295 ;
        RECT 1.615 1.625 2.675 1.665 ;
        RECT 0.095 1.495 2.675 1.625 ;
        RECT 0.095 1.445 1.840 1.495 ;
        RECT 2.505 0.825 2.675 1.495 ;
        RECT 1.945 0.655 2.675 0.825 ;
        RECT 1.945 0.505 2.125 0.655 ;
        RECT 0.820 0.255 2.125 0.505 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 1.435 2.255 1.810 2.635 ;
        RECT 0.595 2.085 0.825 2.125 ;
        RECT 0.595 2.035 1.210 2.085 ;
        RECT 1.955 2.035 2.125 2.165 ;
        RECT 0.595 1.835 2.125 2.035 ;
        RECT 2.360 1.855 2.625 2.635 ;
        RECT 0.595 1.795 1.475 1.835 ;
        RECT 0.095 0.085 0.545 0.595 ;
        RECT 2.305 0.085 2.635 0.485 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__a22oi_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a22oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.075 3.100 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.390 1.075 4.500 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.070 1.075 1.700 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.150 1.075 0.780 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.395 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.141000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.655 0.345 2.465 ;
        RECT 0.935 1.655 1.265 2.125 ;
        RECT 1.775 1.655 2.160 2.125 ;
        RECT 0.095 1.485 2.160 1.655 ;
        RECT 1.870 0.845 2.160 1.485 ;
        RECT 1.355 0.675 3.045 0.845 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.515 2.295 2.625 2.465 ;
        RECT 0.515 1.825 0.765 2.295 ;
        RECT 1.435 1.825 1.605 2.295 ;
        RECT 2.375 1.655 2.625 2.295 ;
        RECT 2.795 1.825 2.965 2.635 ;
        RECT 3.135 1.655 3.465 2.465 ;
        RECT 3.635 1.825 3.805 2.635 ;
        RECT 3.975 1.655 4.305 2.465 ;
        RECT 2.375 1.485 4.305 1.655 ;
        RECT 0.095 0.680 1.185 0.850 ;
        RECT 0.095 0.255 0.345 0.680 ;
        RECT 0.515 0.085 0.845 0.510 ;
        RECT 1.015 0.505 1.185 0.680 ;
        RECT 3.215 0.680 4.375 0.850 ;
        RECT 3.215 0.505 3.385 0.680 ;
        RECT 1.015 0.255 2.105 0.505 ;
        RECT 2.295 0.255 3.385 0.505 ;
        RECT 3.555 0.085 3.885 0.510 ;
        RECT 4.055 0.255 4.375 0.680 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__a22oi_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a22oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a22oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 4.275 1.075 5.685 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 5.910 1.075 7.735 1.285 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 2.615 1.075 4.040 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 1.895 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.755 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.625 0.805 2.125 ;
        RECT 1.395 1.625 1.645 2.125 ;
        RECT 2.235 1.625 2.485 2.125 ;
        RECT 3.075 1.625 3.325 2.125 ;
        RECT 0.595 1.445 3.325 1.625 ;
        RECT 2.195 0.885 2.445 1.445 ;
        RECT 2.195 0.645 5.565 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.090 2.295 4.265 2.465 ;
        RECT 0.090 1.455 0.425 2.295 ;
        RECT 0.975 1.795 1.225 2.295 ;
        RECT 1.815 1.795 2.065 2.295 ;
        RECT 2.655 1.795 2.905 2.295 ;
        RECT 3.495 1.625 4.265 2.295 ;
        RECT 4.435 1.795 4.685 2.635 ;
        RECT 4.855 1.625 5.105 2.465 ;
        RECT 5.275 1.795 5.525 2.635 ;
        RECT 5.695 1.625 5.945 2.465 ;
        RECT 6.115 1.795 6.365 2.635 ;
        RECT 6.535 1.625 6.785 2.465 ;
        RECT 6.955 1.795 7.205 2.635 ;
        RECT 7.375 1.625 7.625 2.465 ;
        RECT 3.495 1.455 7.625 1.625 ;
        RECT 0.095 0.725 2.025 0.905 ;
        RECT 0.095 0.255 0.425 0.725 ;
        RECT 0.595 0.085 0.765 0.555 ;
        RECT 0.935 0.255 1.265 0.725 ;
        RECT 1.435 0.085 1.605 0.555 ;
        RECT 1.775 0.475 2.025 0.725 ;
        RECT 5.735 0.725 7.665 0.905 ;
        RECT 5.735 0.475 5.985 0.725 ;
        RECT 1.775 0.255 3.785 0.475 ;
        RECT 3.975 0.255 5.985 0.475 ;
        RECT 6.155 0.085 6.325 0.555 ;
        RECT 6.495 0.255 6.825 0.725 ;
        RECT 6.995 0.085 7.165 0.555 ;
        RECT 7.335 0.255 7.665 0.725 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
  END
END sky130_fd_sc_hd__a22oi_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a31o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.895 0.995 2.160 1.655 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.415 0.995 1.700 1.655 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.325 1.240 1.655 ;
        RECT 0.935 0.995 1.240 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.375 0.995 2.620 1.655 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.925 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.437250 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.575 0.425 2.425 ;
        RECT 0.095 0.810 0.285 1.575 ;
        RECT 0.095 0.300 0.425 0.810 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.595 1.495 0.845 2.635 ;
        RECT 1.035 1.995 1.285 2.415 ;
        RECT 1.515 2.165 1.845 2.635 ;
        RECT 2.075 1.995 2.325 2.415 ;
        RECT 1.035 1.825 2.325 1.995 ;
        RECT 2.505 1.995 2.835 2.425 ;
        RECT 2.505 1.825 2.960 1.995 ;
        RECT 0.455 0.995 0.765 1.325 ;
        RECT 0.595 0.825 0.765 0.995 ;
        RECT 2.790 0.825 2.960 1.825 ;
        RECT 0.595 0.655 2.960 0.825 ;
        RECT 0.595 0.085 0.925 0.485 ;
        RECT 1.975 0.315 2.305 0.655 ;
        RECT 2.475 0.085 2.805 0.485 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__a31o_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a31o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.185 0.870 2.355 1.325 ;
        RECT 1.965 0.700 2.355 0.870 ;
        RECT 1.965 0.415 2.175 0.700 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.625 1.245 1.795 1.260 ;
        RECT 1.625 1.075 1.955 1.245 ;
        RECT 1.625 0.865 1.795 1.075 ;
        RECT 1.530 0.695 1.795 0.865 ;
        RECT 1.530 0.400 1.700 0.695 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.995 1.395 1.325 ;
        RECT 1.065 0.760 1.270 0.995 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.895 0.755 3.090 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.215 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.595 2.005 0.765 2.465 ;
        RECT 0.090 1.835 0.765 2.005 ;
        RECT 0.090 0.885 0.345 1.835 ;
        RECT 0.090 0.715 0.765 0.885 ;
        RECT 0.595 0.255 0.765 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.135 2.175 0.385 2.635 ;
        RECT 0.935 1.835 1.185 2.635 ;
        RECT 1.355 2.005 1.605 2.425 ;
        RECT 1.815 2.175 2.145 2.635 ;
        RECT 2.335 2.005 2.585 2.425 ;
        RECT 1.355 1.835 2.645 2.005 ;
        RECT 2.875 1.665 3.045 2.465 ;
        RECT 0.555 1.495 3.045 1.665 ;
        RECT 0.555 1.245 0.725 1.495 ;
        RECT 0.555 1.075 0.885 1.245 ;
        RECT 0.090 0.085 0.345 0.545 ;
        RECT 1.015 0.465 1.185 0.545 ;
        RECT 2.535 0.505 2.705 1.495 ;
        RECT 0.955 0.085 1.285 0.465 ;
        RECT 2.375 0.335 2.705 0.505 ;
        RECT 2.460 0.255 2.705 0.335 ;
        RECT 2.875 0.085 3.135 0.565 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__a31o_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a31o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.075 1.705 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.725 1.075 1.055 1.245 ;
        RECT 1.985 1.075 2.315 1.275 ;
        RECT 0.805 0.905 0.975 1.075 ;
        RECT 1.985 0.905 2.170 1.075 ;
        RECT 0.805 0.735 2.170 0.905 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.150 1.445 2.855 1.615 ;
        RECT 0.150 1.075 0.525 1.445 ;
        RECT 2.525 1.075 2.855 1.445 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.575 1.075 4.030 1.285 ;
        RECT 3.815 0.745 4.030 1.075 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.195 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 4.595 1.955 4.765 2.465 ;
        RECT 5.435 1.955 5.605 2.465 ;
        RECT 4.535 1.785 6.295 1.955 ;
        RECT 6.125 0.825 6.295 1.785 ;
        RECT 4.505 0.655 6.295 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.175 1.955 0.345 2.465 ;
        RECT 0.515 2.125 0.845 2.635 ;
        RECT 1.015 1.955 1.185 2.465 ;
        RECT 1.355 2.125 1.685 2.635 ;
        RECT 1.855 1.955 2.025 2.465 ;
        RECT 2.195 2.125 2.525 2.635 ;
        RECT 2.815 2.295 3.825 2.465 ;
        RECT 2.815 1.955 2.985 2.295 ;
        RECT 0.175 1.785 2.985 1.955 ;
        RECT 3.155 1.625 3.485 2.115 ;
        RECT 3.655 1.795 3.825 2.295 ;
        RECT 4.095 2.125 4.425 2.635 ;
        RECT 4.935 2.125 5.265 2.635 ;
        RECT 5.775 2.125 6.105 2.635 ;
        RECT 3.155 1.455 4.395 1.625 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 3.155 0.870 3.345 1.455 ;
        RECT 4.225 1.325 4.395 1.455 ;
        RECT 4.225 0.995 5.935 1.325 ;
        RECT 2.350 0.805 3.345 0.870 ;
        RECT 2.350 0.700 3.485 0.805 ;
        RECT 2.350 0.565 2.520 0.700 ;
        RECT 1.355 0.395 2.520 0.565 ;
        RECT 2.700 0.085 2.985 0.530 ;
        RECT 3.155 0.295 3.485 0.700 ;
        RECT 3.735 0.085 4.265 0.565 ;
        RECT 4.935 0.085 5.265 0.485 ;
        RECT 5.775 0.085 6.105 0.485 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
END sky130_fd_sc_hd__a31o_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a31oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.070 1.445 1.455 1.665 ;
        RECT 1.270 0.995 1.455 1.445 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.610 0.335 1.055 1.275 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.365 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.965 0.995 2.215 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.295 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.481250 ;
    PORT
      LAYER li1 ;
        RECT 1.875 1.665 2.210 2.445 ;
        RECT 1.625 1.495 2.210 1.665 ;
        RECT 1.625 0.825 1.795 1.495 ;
        RECT 1.380 0.715 1.795 0.825 ;
        RECT 1.380 0.295 1.785 0.715 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.090 1.495 0.420 2.635 ;
        RECT 0.590 2.005 0.765 2.415 ;
        RECT 0.935 2.175 1.265 2.635 ;
        RECT 1.470 2.005 1.695 2.415 ;
        RECT 0.590 1.835 1.695 2.005 ;
        RECT 0.090 0.085 0.430 0.815 ;
        RECT 1.955 0.085 2.215 0.565 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__a31oi_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a31oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.955 0.995 2.665 1.615 ;
        RECT 2.905 0.995 3.075 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.050 0.995 1.755 1.615 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.995 0.820 1.615 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.265 1.275 4.490 1.625 ;
        RECT 3.820 1.075 4.490 1.275 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.595 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.922000 ;
    PORT
      LAYER li1 ;
        RECT 3.755 1.615 4.085 2.115 ;
        RECT 3.255 1.445 4.085 1.615 ;
        RECT 3.255 0.825 3.570 1.445 ;
        RECT 2.295 0.655 4.505 0.825 ;
        RECT 3.255 0.255 3.425 0.655 ;
        RECT 4.175 0.295 4.505 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.175 1.955 0.345 2.465 ;
        RECT 0.515 2.125 0.845 2.635 ;
        RECT 1.015 1.955 1.185 2.465 ;
        RECT 1.355 2.125 1.685 2.635 ;
        RECT 1.855 1.955 2.025 2.465 ;
        RECT 2.310 2.125 2.980 2.635 ;
        RECT 3.335 2.295 4.425 2.465 ;
        RECT 3.335 1.955 3.505 2.295 ;
        RECT 0.175 1.785 3.505 1.955 ;
        RECT 4.255 1.795 4.425 2.295 ;
        RECT 0.095 0.655 2.105 0.825 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.355 0.295 3.075 0.465 ;
        RECT 3.675 0.085 4.005 0.465 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__a31oi_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a31oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a31oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.825 0.995 5.420 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.995 3.550 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.120 0.995 1.735 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 5.670 0.995 6.855 1.630 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.815 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.443500 ;
    PORT
      LAYER li1 ;
        RECT 6.075 1.915 7.245 2.085 ;
        RECT 7.045 0.805 7.245 1.915 ;
        RECT 3.975 0.635 7.585 0.805 ;
        RECT 6.575 0.255 6.745 0.635 ;
        RECT 7.415 0.255 7.585 0.635 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.175 1.665 0.345 2.465 ;
        RECT 0.515 1.915 0.845 2.635 ;
        RECT 1.015 1.665 1.185 2.465 ;
        RECT 1.355 1.915 1.685 2.635 ;
        RECT 1.855 1.665 2.025 2.465 ;
        RECT 2.195 1.915 2.525 2.635 ;
        RECT 2.695 1.665 2.865 2.465 ;
        RECT 3.035 1.915 3.365 2.635 ;
        RECT 3.535 1.665 3.705 2.465 ;
        RECT 3.895 1.915 4.225 2.635 ;
        RECT 4.395 1.665 4.565 2.465 ;
        RECT 4.735 2.255 5.065 2.635 ;
        RECT 5.235 2.425 5.405 2.465 ;
        RECT 5.235 2.255 7.665 2.425 ;
        RECT 5.235 1.665 5.405 2.255 ;
        RECT 0.175 1.495 5.405 1.665 ;
        RECT 7.415 1.495 7.665 2.255 ;
        RECT 0.175 0.635 3.785 0.805 ;
        RECT 0.175 0.255 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.255 1.185 0.635 ;
        RECT 1.355 0.085 1.685 0.465 ;
        RECT 1.855 0.255 2.025 0.635 ;
        RECT 2.195 0.295 5.565 0.465 ;
        RECT 6.075 0.085 6.405 0.465 ;
        RECT 6.915 0.085 7.245 0.465 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
  END
END sky130_fd_sc_hd__a31oi_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a32o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.990 0.665 2.280 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.530 0.665 1.800 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.070 0.995 1.320 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.450 0.660 2.870 1.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.325 1.325 3.530 1.615 ;
        RECT 3.180 0.995 3.530 1.325 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.675 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.544500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.915 0.425 2.425 ;
        RECT 0.090 0.560 0.345 1.915 ;
        RECT 0.090 0.300 0.425 0.560 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.675 1.835 1.005 2.635 ;
        RECT 1.250 2.045 1.535 2.465 ;
        RECT 1.790 2.215 2.120 2.635 ;
        RECT 2.345 2.295 3.505 2.465 ;
        RECT 2.345 2.045 2.675 2.295 ;
        RECT 1.250 1.875 2.675 2.045 ;
        RECT 2.905 1.665 3.075 2.125 ;
        RECT 3.335 1.795 3.505 2.295 ;
        RECT 0.705 1.495 3.075 1.665 ;
        RECT 0.705 1.325 0.875 1.495 ;
        RECT 0.570 0.995 0.875 1.325 ;
        RECT 0.705 0.825 0.875 0.995 ;
        RECT 0.705 0.655 1.265 0.825 ;
        RECT 1.095 0.485 1.265 0.655 ;
        RECT 0.595 0.085 0.925 0.485 ;
        RECT 1.095 0.315 2.710 0.485 ;
        RECT 3.255 0.085 3.585 0.805 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__a32o_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a32o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.685 0.955 2.985 1.325 ;
        RECT 2.755 0.610 2.985 0.955 ;
        RECT 2.755 0.415 3.105 0.610 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.305 1.325 3.545 1.625 ;
        RECT 3.165 0.995 3.545 1.325 ;
        RECT 3.305 0.425 3.545 0.995 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.815 0.995 4.055 1.630 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.345 1.445 2.550 1.615 ;
        RECT 2.345 1.245 2.515 1.445 ;
        RECT 2.085 1.075 2.515 1.245 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.115 0.745 1.530 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.135 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.695500 ;
    PORT
      LAYER li1 ;
        RECT 0.135 1.955 0.345 2.465 ;
        RECT 1.015 1.955 1.185 2.465 ;
        RECT 0.135 1.785 1.185 1.955 ;
        RECT 0.135 0.825 0.345 1.785 ;
        RECT 0.135 0.655 0.845 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.515 2.125 0.845 2.635 ;
        RECT 1.535 2.295 2.545 2.465 ;
        RECT 1.535 1.785 1.705 2.295 ;
        RECT 1.875 1.945 2.205 2.115 ;
        RECT 2.375 1.965 2.545 2.295 ;
        RECT 2.715 2.140 3.045 2.635 ;
        RECT 3.375 1.965 3.545 2.465 ;
        RECT 1.875 1.615 2.125 1.945 ;
        RECT 2.375 1.795 3.545 1.965 ;
        RECT 3.715 1.915 4.050 2.635 ;
        RECT 0.535 1.445 2.125 1.615 ;
        RECT 0.535 0.995 0.705 1.445 ;
        RECT 1.700 0.785 1.890 1.445 ;
        RECT 1.700 0.615 2.585 0.785 ;
        RECT 0.090 0.085 0.425 0.465 ;
        RECT 0.935 0.085 1.640 0.445 ;
        RECT 2.255 0.275 2.585 0.615 ;
        RECT 3.715 0.085 4.050 0.805 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__a32o_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a32o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.280 1.075 5.075 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.335 1.075 4.030 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.210 1.075 3.105 1.295 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 5.630 1.075 6.780 1.625 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 7.030 1.295 7.225 1.635 ;
        RECT 7.030 1.075 7.710 1.295 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.815 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.665 0.765 2.465 ;
        RECT 1.435 1.665 1.605 2.465 ;
        RECT 0.120 1.495 1.605 1.665 ;
        RECT 0.120 0.805 0.340 1.495 ;
        RECT 0.120 0.635 1.605 0.805 ;
        RECT 0.595 0.255 0.765 0.635 ;
        RECT 1.435 0.255 1.605 0.635 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.095 1.915 0.425 2.635 ;
        RECT 0.935 1.915 1.265 2.635 ;
        RECT 1.775 1.915 2.105 2.635 ;
        RECT 2.275 2.085 2.445 2.465 ;
        RECT 2.615 2.255 2.945 2.635 ;
        RECT 3.215 2.085 3.385 2.465 ;
        RECT 3.555 2.255 3.885 2.635 ;
        RECT 4.055 2.085 4.225 2.465 ;
        RECT 4.395 2.255 4.725 2.635 ;
        RECT 4.895 2.255 7.725 2.425 ;
        RECT 4.895 2.085 5.065 2.255 ;
        RECT 2.275 1.915 5.065 2.085 ;
        RECT 6.135 2.075 7.305 2.085 ;
        RECT 5.280 1.915 7.305 2.075 ;
        RECT 5.280 1.905 6.200 1.915 ;
        RECT 5.280 1.665 5.450 1.905 ;
        RECT 7.475 1.755 7.725 2.255 ;
        RECT 1.800 1.495 5.450 1.665 ;
        RECT 1.800 1.325 1.970 1.495 ;
        RECT 0.570 0.995 1.970 1.325 ;
        RECT 2.275 0.655 3.885 0.825 ;
        RECT 5.280 0.805 5.450 1.495 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 1.775 0.085 2.105 0.465 ;
        RECT 2.275 0.255 2.445 0.655 ;
        RECT 4.395 0.635 6.425 0.805 ;
        RECT 6.635 0.645 7.645 0.815 ;
        RECT 6.635 0.465 6.805 0.645 ;
        RECT 2.615 0.085 2.945 0.465 ;
        RECT 3.135 0.295 5.145 0.465 ;
        RECT 5.670 0.295 6.805 0.465 ;
        RECT 6.635 0.255 6.805 0.295 ;
        RECT 6.975 0.085 7.305 0.465 ;
        RECT 7.475 0.255 7.645 0.645 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
  END
END sky130_fd_sc_hd__a32o_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a32oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.230 1.075 1.595 1.255 ;
        RECT 1.405 0.765 1.595 1.075 ;
        RECT 1.405 0.345 1.705 0.765 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.805 0.995 2.165 1.325 ;
        RECT 1.965 0.415 2.165 0.995 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.335 1.015 2.750 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.855 1.425 1.255 1.615 ;
        RECT 0.855 0.995 1.025 1.425 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.345 1.325 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.785 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.575500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.785 0.865 2.085 ;
        RECT 0.515 0.805 0.685 1.785 ;
        RECT 0.515 0.635 1.165 0.805 ;
        RECT 0.915 0.295 1.165 0.635 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 2.255 1.345 2.465 ;
        RECT 0.085 1.835 0.345 2.255 ;
        RECT 1.095 1.955 1.345 2.255 ;
        RECT 1.555 2.135 1.805 2.635 ;
        RECT 2.015 1.955 2.185 2.465 ;
        RECT 1.095 1.785 2.185 1.955 ;
        RECT 2.015 1.745 2.185 1.785 ;
        RECT 2.355 1.495 2.695 2.635 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 2.355 0.085 2.695 0.805 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__a32oi_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a32oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.415 1.075 3.220 1.625 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.725 1.075 4.480 1.625 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.715 1.075 5.860 1.625 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.080 1.725 1.285 ;
        RECT 1.175 1.075 1.505 1.080 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 1.285 0.325 1.625 ;
        RECT 0.145 1.075 0.825 1.285 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.975 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.955 0.845 2.125 ;
        RECT 0.595 1.625 0.765 1.955 ;
        RECT 1.435 1.625 1.605 2.125 ;
        RECT 0.595 1.455 2.180 1.625 ;
        RECT 1.965 0.825 2.180 1.455 ;
        RECT 1.355 0.655 3.100 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.175 2.295 2.025 2.465 ;
        RECT 0.175 1.795 0.345 2.295 ;
        RECT 1.015 1.795 1.185 2.295 ;
        RECT 1.855 2.085 2.025 2.295 ;
        RECT 2.270 2.255 2.940 2.635 ;
        RECT 3.180 2.085 3.350 2.465 ;
        RECT 3.550 2.255 4.220 2.635 ;
        RECT 4.390 2.085 4.560 2.465 ;
        RECT 4.765 2.255 5.435 2.635 ;
        RECT 5.635 2.085 5.805 2.465 ;
        RECT 1.855 1.915 5.805 2.085 ;
        RECT 1.855 1.795 2.025 1.915 ;
        RECT 3.180 1.795 3.350 1.915 ;
        RECT 4.390 1.795 4.560 1.915 ;
        RECT 5.635 1.795 5.805 1.915 ;
        RECT 0.175 0.715 1.185 0.885 ;
        RECT 0.175 0.465 0.345 0.715 ;
        RECT 0.095 0.295 0.425 0.465 ;
        RECT 0.595 0.085 0.765 0.545 ;
        RECT 1.015 0.465 1.185 0.715 ;
        RECT 3.620 0.635 5.390 0.805 ;
        RECT 0.935 0.295 2.115 0.465 ;
        RECT 2.350 0.295 4.370 0.465 ;
        RECT 4.555 0.085 4.890 0.465 ;
        RECT 5.060 0.275 5.390 0.635 ;
        RECT 5.560 0.085 5.885 0.885 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
END sky130_fd_sc_hd__a32oi_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a32oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a32oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.775 1.075 5.465 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.095 1.075 7.695 1.300 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 8.295 1.075 9.985 1.280 ;
        RECT 9.805 0.755 9.985 1.075 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 2.585 0.995 3.555 1.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.305 0.330 1.965 ;
        RECT 0.110 1.075 1.750 1.305 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 10.115 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.745 0.845 2.085 ;
        RECT 1.355 1.745 1.685 2.085 ;
        RECT 1.975 1.745 2.525 2.085 ;
        RECT 3.035 1.745 3.365 2.085 ;
        RECT 0.515 1.575 3.365 1.745 ;
        RECT 1.975 0.990 2.365 1.575 ;
        RECT 2.195 0.805 2.365 0.990 ;
        RECT 2.195 0.635 5.565 0.805 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.095 2.255 3.705 2.425 ;
        RECT 3.535 1.745 3.705 2.255 ;
        RECT 3.895 1.915 4.225 2.635 ;
        RECT 4.395 1.745 4.565 2.465 ;
        RECT 4.770 1.915 5.440 2.635 ;
        RECT 5.640 1.745 5.810 2.465 ;
        RECT 6.215 1.915 6.545 2.635 ;
        RECT 6.715 1.745 6.885 2.465 ;
        RECT 7.055 1.915 7.385 2.635 ;
        RECT 7.555 1.745 7.725 2.465 ;
        RECT 8.415 1.915 8.745 2.635 ;
        RECT 8.915 1.745 9.085 2.465 ;
        RECT 9.255 1.915 9.585 2.635 ;
        RECT 9.755 1.745 9.925 2.465 ;
        RECT 3.535 1.575 9.925 1.745 ;
        RECT 0.175 0.635 2.025 0.805 ;
        RECT 6.215 0.635 9.505 0.805 ;
        RECT 0.175 0.255 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.255 1.185 0.635 ;
        RECT 1.855 0.465 2.025 0.635 ;
        RECT 1.355 0.085 1.685 0.465 ;
        RECT 1.855 0.295 3.785 0.465 ;
        RECT 3.975 0.295 7.805 0.465 ;
        RECT 7.995 0.085 8.325 0.465 ;
        RECT 8.495 0.255 8.665 0.635 ;
        RECT 8.835 0.085 9.165 0.465 ;
        RECT 9.335 0.255 9.505 0.635 ;
        RECT 9.685 0.085 10.025 0.465 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
  END
END sky130_fd_sc_hd__a32oi_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a41o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.535 1.325 1.835 1.620 ;
        RECT 1.535 0.995 1.915 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.225 0.600 2.445 1.325 ;
        RECT 1.700 0.415 2.650 0.600 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.705 0.995 3.085 1.625 ;
        RECT 2.880 0.395 3.085 0.995 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.315 0.995 3.570 1.625 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.075 1.335 1.635 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.675 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.165 0.425 2.425 ;
        RECT 0.085 0.560 0.345 2.165 ;
        RECT 0.085 0.300 0.425 0.560 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.595 2.175 0.845 2.635 ;
        RECT 1.035 1.995 1.365 2.425 ;
        RECT 0.515 1.825 1.365 1.995 ;
        RECT 1.535 1.965 1.705 2.465 ;
        RECT 1.915 2.175 2.165 2.635 ;
        RECT 2.375 1.965 2.545 2.465 ;
        RECT 2.845 2.175 3.095 2.635 ;
        RECT 3.335 1.965 3.505 2.465 ;
        RECT 0.515 0.905 0.685 1.825 ;
        RECT 1.535 1.795 3.505 1.965 ;
        RECT 0.515 0.810 1.335 0.905 ;
        RECT 0.515 0.735 1.530 0.810 ;
        RECT 0.595 0.085 0.925 0.565 ;
        RECT 1.115 0.300 1.530 0.735 ;
        RECT 3.255 0.085 3.595 0.810 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__a41o_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a41o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.785 0.730 4.005 1.625 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.335 1.245 3.550 1.625 ;
        RECT 3.085 1.075 3.550 1.245 ;
        RECT 3.335 0.745 3.550 1.075 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.685 1.435 3.090 1.625 ;
        RECT 2.685 0.995 2.855 1.435 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.000 0.995 2.335 1.625 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.400 1.075 1.730 1.295 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.135 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.755 0.785 2.465 ;
        RECT 0.595 0.295 0.765 0.755 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.095 1.495 0.425 2.635 ;
        RECT 1.015 1.835 1.265 2.635 ;
        RECT 1.455 1.665 1.785 2.425 ;
        RECT 1.955 1.965 2.125 2.465 ;
        RECT 2.335 2.175 2.585 2.635 ;
        RECT 2.795 1.965 2.965 2.465 ;
        RECT 3.335 2.175 3.585 2.635 ;
        RECT 3.795 1.965 3.965 2.465 ;
        RECT 1.955 1.795 3.965 1.965 ;
        RECT 0.980 1.495 1.785 1.665 ;
        RECT 0.980 0.805 1.150 1.495 ;
        RECT 0.095 0.085 0.425 0.805 ;
        RECT 0.980 0.635 2.545 0.805 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 1.495 0.255 1.705 0.635 ;
        RECT 2.375 0.465 2.545 0.635 ;
        RECT 1.875 0.085 2.205 0.465 ;
        RECT 2.375 0.295 4.045 0.465 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__a41o_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a41o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.075 4.065 1.295 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.275 1.075 4.975 1.285 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 5.155 1.075 6.185 1.295 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 6.495 1.075 7.505 1.295 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.075 3.145 1.280 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.455 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.745 0.765 2.465 ;
        RECT 1.435 1.745 1.605 2.465 ;
        RECT 0.150 1.575 1.605 1.745 ;
        RECT 0.150 0.805 0.320 1.575 ;
        RECT 0.150 0.635 1.605 0.805 ;
        RECT 0.595 0.255 0.765 0.635 ;
        RECT 1.435 0.255 1.605 0.635 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.095 1.915 0.425 2.635 ;
        RECT 0.935 1.915 1.265 2.635 ;
        RECT 1.775 1.915 2.125 2.635 ;
        RECT 2.375 2.295 3.405 2.465 ;
        RECT 2.375 1.795 2.545 2.295 ;
        RECT 2.715 1.955 3.045 2.125 ;
        RECT 2.795 1.625 2.965 1.955 ;
        RECT 1.775 1.455 2.965 1.625 ;
        RECT 3.235 1.705 3.405 2.295 ;
        RECT 3.575 1.915 3.905 2.635 ;
        RECT 4.075 1.705 4.245 2.465 ;
        RECT 4.415 1.915 4.745 2.635 ;
        RECT 4.935 1.705 5.105 2.465 ;
        RECT 5.345 1.915 6.035 2.635 ;
        RECT 6.275 1.705 6.445 2.465 ;
        RECT 6.615 1.915 6.945 2.635 ;
        RECT 7.115 1.705 7.285 2.465 ;
        RECT 3.235 1.535 7.370 1.705 ;
        RECT 1.775 1.245 1.945 1.455 ;
        RECT 0.490 1.075 1.945 1.245 ;
        RECT 1.775 0.815 1.945 1.075 ;
        RECT 1.775 0.645 3.905 0.815 ;
        RECT 4.075 0.645 5.165 0.815 ;
        RECT 5.355 0.645 7.285 0.815 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 1.775 0.085 2.125 0.465 ;
        RECT 2.295 0.255 2.465 0.645 ;
        RECT 4.075 0.465 4.245 0.645 ;
        RECT 2.635 0.085 2.965 0.465 ;
        RECT 3.155 0.295 4.245 0.465 ;
        RECT 4.415 0.295 6.105 0.465 ;
        RECT 6.615 0.085 6.945 0.465 ;
        RECT 7.115 0.255 7.285 0.645 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
  END
END sky130_fd_sc_hd__a41o_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a41oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.780 0.995 3.085 1.615 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.890 0.755 2.210 1.665 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.470 0.755 1.710 1.665 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.960 0.965 1.250 1.665 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.540 0.965 0.780 1.665 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.215 1.015 ;
        RECT 0.150 0.065 1.060 0.105 ;
        RECT 0.150 -0.085 0.320 0.065 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.669500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.845 0.425 2.425 ;
        RECT 0.090 0.785 0.360 1.845 ;
        RECT 0.090 0.615 1.290 0.785 ;
        RECT 0.090 0.285 0.345 0.615 ;
        RECT 1.120 0.465 1.290 0.615 ;
        RECT 2.685 0.465 3.015 0.805 ;
        RECT 1.120 0.295 3.015 0.465 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.595 2.015 0.845 2.465 ;
        RECT 1.120 2.195 1.450 2.635 ;
        RECT 1.760 2.015 1.930 2.465 ;
        RECT 2.215 2.195 2.545 2.635 ;
        RECT 2.765 2.015 3.015 2.465 ;
        RECT 0.595 1.845 3.015 2.015 ;
        RECT 0.620 0.085 0.950 0.445 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__a41oi_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a41oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.785 1.075 2.455 1.295 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.665 1.075 3.365 1.285 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.545 1.075 4.575 1.295 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.755 1.075 5.895 1.295 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.075 1.555 1.280 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.095 0.105 5.845 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.621000 ;
    PORT
      LAYER li1 ;
        RECT 1.125 1.625 1.455 2.125 ;
        RECT 0.145 1.455 1.455 1.625 ;
        RECT 0.145 0.815 0.315 1.455 ;
        RECT 0.145 0.645 2.295 0.815 ;
        RECT 0.685 0.255 0.855 0.645 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.785 2.295 1.795 2.465 ;
        RECT 0.785 1.795 0.955 2.295 ;
        RECT 1.625 1.705 1.795 2.295 ;
        RECT 1.965 1.915 2.295 2.635 ;
        RECT 2.465 1.705 2.635 2.465 ;
        RECT 2.805 1.915 3.135 2.635 ;
        RECT 3.325 1.705 3.495 2.465 ;
        RECT 3.755 1.915 4.425 2.635 ;
        RECT 4.665 1.705 4.835 2.465 ;
        RECT 5.005 1.915 5.335 2.635 ;
        RECT 5.505 1.705 5.675 2.465 ;
        RECT 1.625 1.535 5.760 1.705 ;
        RECT 2.465 0.645 3.555 0.815 ;
        RECT 3.745 0.645 5.675 0.815 ;
        RECT 2.465 0.465 2.635 0.645 ;
        RECT 0.185 0.085 0.515 0.465 ;
        RECT 1.025 0.085 1.375 0.465 ;
        RECT 1.545 0.295 2.635 0.465 ;
        RECT 2.805 0.295 4.495 0.465 ;
        RECT 5.005 0.085 5.335 0.465 ;
        RECT 5.505 0.255 5.675 0.645 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
END sky130_fd_sc_hd__a41oi_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a41oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a41oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 2.385 0.995 4.205 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 4.405 1.075 6.315 1.285 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.560 1.075 7.955 1.300 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 8.285 1.075 9.975 1.280 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.305 0.325 1.965 ;
        RECT 0.105 1.075 1.745 1.305 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 10.115 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.745 0.845 2.085 ;
        RECT 1.350 1.745 1.685 2.085 ;
        RECT 0.515 1.685 1.685 1.745 ;
        RECT 0.515 1.575 2.155 1.685 ;
        RECT 1.350 1.495 2.155 1.575 ;
        RECT 1.935 0.805 2.155 1.495 ;
        RECT 0.595 0.635 4.015 0.805 ;
        RECT 0.595 0.255 0.765 0.635 ;
        RECT 1.435 0.255 1.605 0.635 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 2.165 2.425 2.335 2.465 ;
        RECT 0.090 2.255 2.335 2.425 ;
        RECT 2.505 2.255 3.175 2.635 ;
        RECT 2.165 2.075 2.335 2.255 ;
        RECT 3.345 2.075 3.515 2.465 ;
        RECT 2.165 1.905 3.515 2.075 ;
        RECT 3.685 1.915 4.015 2.635 ;
        RECT 3.345 1.745 3.515 1.905 ;
        RECT 4.185 1.745 4.355 2.425 ;
        RECT 4.620 1.915 4.950 2.635 ;
        RECT 5.120 1.745 5.290 2.465 ;
        RECT 5.495 1.915 6.165 2.635 ;
        RECT 6.385 1.745 6.555 2.465 ;
        RECT 6.725 1.915 7.055 2.635 ;
        RECT 7.225 1.745 7.395 2.465 ;
        RECT 7.565 1.915 7.895 2.635 ;
        RECT 8.065 1.745 8.235 2.465 ;
        RECT 8.405 1.915 8.735 2.635 ;
        RECT 8.905 1.745 9.075 2.465 ;
        RECT 9.245 1.915 9.575 2.635 ;
        RECT 9.775 1.745 9.945 2.465 ;
        RECT 3.345 1.575 9.945 1.745 ;
        RECT 4.525 0.635 7.895 0.805 ;
        RECT 8.065 0.635 9.915 0.805 ;
        RECT 8.065 0.465 8.235 0.635 ;
        RECT 0.090 0.085 0.425 0.465 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 1.775 0.085 2.105 0.465 ;
        RECT 2.425 0.295 6.115 0.465 ;
        RECT 6.305 0.295 8.235 0.465 ;
        RECT 8.065 0.255 8.235 0.295 ;
        RECT 8.405 0.085 8.735 0.465 ;
        RECT 8.905 0.255 9.075 0.635 ;
        RECT 9.245 0.085 9.575 0.465 ;
        RECT 9.745 0.255 9.915 0.635 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
  END
END sky130_fd_sc_hd__a41oi_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a211o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.485 0.995 2.060 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.025 0.995 1.305 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.240 0.995 2.675 1.325 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.855 0.995 3.125 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.215 1.015 ;
        RECT 0.135 -0.085 0.305 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.437250 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.685 0.355 2.455 ;
        RECT 0.090 0.265 0.425 1.685 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.525 1.915 0.855 2.635 ;
        RECT 1.045 2.095 1.305 2.455 ;
        RECT 1.475 2.265 1.805 2.635 ;
        RECT 1.975 2.095 2.235 2.455 ;
        RECT 1.045 1.865 2.235 2.095 ;
        RECT 2.805 1.685 3.095 2.455 ;
        RECT 0.600 1.505 3.095 1.685 ;
        RECT 0.600 0.815 0.825 1.505 ;
        RECT 0.600 0.625 3.085 0.815 ;
        RECT 0.605 0.085 1.350 0.455 ;
        RECT 1.915 0.265 2.170 0.625 ;
        RECT 2.350 0.085 2.680 0.455 ;
        RECT 2.860 0.265 3.085 0.625 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__a211o_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a211o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.980 1.045 2.450 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.480 1.045 1.810 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.620 1.045 3.070 1.275 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.260 1.045 3.595 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.675 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.452000 ;
    PORT
      LAYER li1 ;
        RECT 0.555 0.635 0.785 2.335 ;
        RECT 0.555 0.255 0.775 0.635 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.090 1.490 0.385 2.635 ;
        RECT 1.000 1.830 1.255 2.635 ;
        RECT 1.455 2.020 1.785 2.465 ;
        RECT 1.955 2.190 2.230 2.635 ;
        RECT 2.465 2.020 2.795 2.465 ;
        RECT 1.455 1.840 2.795 2.020 ;
        RECT 3.255 1.660 3.585 2.325 ;
        RECT 1.000 1.490 3.585 1.660 ;
        RECT 0.090 0.085 0.385 0.905 ;
        RECT 1.000 0.875 1.310 1.490 ;
        RECT 1.000 0.695 3.585 0.875 ;
        RECT 0.945 0.085 1.795 0.445 ;
        RECT 2.275 0.275 2.605 0.695 ;
        RECT 2.810 0.085 3.085 0.525 ;
        RECT 3.255 0.275 3.585 0.695 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__a211o_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a211o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 5.035 1.020 5.380 1.330 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.495 1.510 5.845 1.700 ;
        RECT 4.495 1.020 4.825 1.510 ;
        RECT 5.635 1.320 5.845 1.510 ;
        RECT 5.635 1.020 6.225 1.320 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.625 1.445 4.175 1.700 ;
        RECT 2.625 1.325 2.805 1.445 ;
        RECT 2.540 0.985 2.805 1.325 ;
        RECT 3.845 0.985 4.175 1.445 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.975 0.985 3.645 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.933750 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.705 0.780 2.465 ;
        RECT 1.450 1.705 1.640 2.465 ;
        RECT 0.085 1.495 1.640 1.705 ;
        RECT 0.085 0.875 0.340 1.495 ;
        RECT 0.085 0.635 2.025 0.875 ;
        RECT 0.985 0.615 2.025 0.635 ;
        RECT 0.985 0.255 1.175 0.615 ;
        RECT 1.845 0.255 2.025 0.615 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 0.395 0.105 6.435 1.015 ;
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.090 1.875 0.425 2.635 ;
        RECT 0.950 1.875 1.280 2.635 ;
        RECT 1.810 1.835 2.060 2.635 ;
        RECT 2.320 2.210 4.450 2.465 ;
        RECT 4.620 2.275 4.950 2.635 ;
        RECT 4.120 2.105 4.450 2.210 ;
        RECT 5.160 2.105 5.420 2.465 ;
        RECT 5.590 2.275 5.920 2.635 ;
        RECT 6.090 2.105 6.345 2.465 ;
        RECT 2.280 1.870 3.510 2.040 ;
        RECT 4.120 1.880 6.345 2.105 ;
        RECT 2.280 1.675 2.455 1.870 ;
        RECT 2.185 1.505 2.455 1.675 ;
        RECT 6.015 1.535 6.345 1.880 ;
        RECT 2.185 1.325 2.370 1.505 ;
        RECT 0.525 1.045 2.370 1.325 ;
        RECT 2.195 0.805 2.370 1.045 ;
        RECT 2.195 0.615 5.490 0.805 ;
        RECT 0.485 0.085 0.815 0.465 ;
        RECT 1.345 0.085 1.675 0.445 ;
        RECT 2.220 0.085 2.555 0.445 ;
        RECT 2.725 0.255 2.970 0.615 ;
        RECT 3.140 0.085 3.470 0.445 ;
        RECT 3.640 0.255 4.020 0.615 ;
        RECT 4.190 0.085 4.560 0.445 ;
        RECT 5.160 0.275 5.490 0.615 ;
        RECT 6.015 0.085 6.345 0.805 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
END sky130_fd_sc_hd__a211o_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a211oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.995 1.245 1.325 ;
        RECT 0.605 0.265 0.855 0.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.765 0.435 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.325 1.755 2.455 ;
        RECT 1.425 0.995 1.755 1.325 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.995 2.235 1.615 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.410 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.619250 ;
    PORT
      LAYER li1 ;
        RECT 1.935 1.785 2.660 2.455 ;
        RECT 2.445 0.815 2.660 1.785 ;
        RECT 1.180 0.625 2.660 0.815 ;
        RECT 1.180 0.265 1.365 0.625 ;
        RECT 2.055 0.265 2.280 0.625 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.250 1.725 0.500 2.455 ;
        RECT 0.670 1.905 1.000 2.635 ;
        RECT 1.170 1.725 1.355 2.455 ;
        RECT 0.250 1.525 1.355 1.725 ;
        RECT 0.085 0.085 0.425 0.595 ;
        RECT 1.545 0.085 1.875 0.455 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__a211oi_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a211oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.370 1.035 3.080 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.175 1.285 4.500 1.655 ;
        RECT 3.740 1.035 4.500 1.285 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.035 1.285 1.255 1.615 ;
        RECT 1.035 1.035 1.785 1.285 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 0.995 0.405 1.615 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.055 0.105 4.525 1.015 ;
        RECT 0.125 -0.085 0.295 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.826000 ;
    PORT
      LAYER li1 ;
        RECT 0.575 1.785 0.905 2.105 ;
        RECT 0.575 0.855 0.855 1.785 ;
        RECT 0.575 0.655 3.145 0.855 ;
        RECT 0.575 0.255 0.835 0.655 ;
        RECT 1.505 0.285 1.695 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.145 2.285 2.215 2.455 ;
        RECT 0.145 1.785 0.405 2.285 ;
        RECT 1.075 2.255 2.215 2.285 ;
        RECT 1.075 1.785 1.265 2.255 ;
        RECT 1.435 1.655 1.765 2.075 ;
        RECT 1.935 1.835 2.215 2.255 ;
        RECT 2.435 1.835 2.665 2.635 ;
        RECT 2.845 1.655 3.115 2.465 ;
        RECT 3.295 1.835 3.525 2.635 ;
        RECT 3.705 1.655 3.975 2.465 ;
        RECT 4.155 1.835 4.385 2.635 ;
        RECT 1.435 1.455 3.975 1.655 ;
        RECT 0.145 0.085 0.395 0.815 ;
        RECT 3.325 0.635 4.435 0.855 ;
        RECT 3.325 0.475 3.495 0.635 ;
        RECT 1.005 0.085 1.335 0.475 ;
        RECT 1.865 0.085 2.195 0.475 ;
        RECT 2.385 0.265 3.495 0.475 ;
        RECT 3.675 0.085 4.005 0.455 ;
        RECT 4.185 0.265 4.435 0.635 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__a211oi_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a211oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a211oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.660 1.245 3.005 1.275 ;
        RECT 1.655 1.075 3.005 1.245 ;
        RECT 1.660 1.035 3.005 1.075 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.445 3.575 1.625 ;
        RECT 0.100 1.035 1.385 1.445 ;
        RECT 3.245 1.035 3.575 1.445 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met1 ;
        RECT 3.770 1.600 4.060 1.645 ;
        RECT 6.530 1.600 6.820 1.645 ;
        RECT 3.770 1.460 6.820 1.600 ;
        RECT 3.770 1.415 4.060 1.460 ;
        RECT 6.530 1.415 6.820 1.460 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.130 1.275 6.350 1.695 ;
        RECT 5.000 1.035 6.350 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.355 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.685000 ;
    PORT
      LAYER li1 ;
        RECT 5.170 1.865 7.275 2.085 ;
        RECT 6.930 1.495 7.275 1.865 ;
        RECT 1.775 0.825 6.355 0.865 ;
        RECT 7.105 0.825 7.275 1.495 ;
        RECT 1.775 0.695 7.275 0.825 ;
        RECT 1.775 0.675 3.330 0.695 ;
        RECT 3.875 0.625 7.275 0.695 ;
        RECT 3.875 0.615 5.045 0.625 ;
        RECT 3.875 0.255 4.195 0.615 ;
        RECT 4.875 0.255 5.045 0.615 ;
        RECT 5.715 0.615 7.275 0.625 ;
        RECT 5.715 0.255 5.885 0.615 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.095 2.085 0.345 2.465 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.015 2.105 1.185 2.465 ;
        RECT 1.355 2.275 1.685 2.635 ;
        RECT 1.855 2.105 2.025 2.465 ;
        RECT 2.195 2.275 2.525 2.635 ;
        RECT 2.695 2.105 2.865 2.465 ;
        RECT 3.035 2.275 3.365 2.635 ;
        RECT 3.535 2.255 7.270 2.465 ;
        RECT 3.535 2.105 3.705 2.255 ;
        RECT 1.015 2.085 3.705 2.105 ;
        RECT 0.095 1.795 3.705 2.085 ;
        RECT 3.875 1.785 4.910 2.085 ;
        RECT 4.630 1.695 4.910 1.785 ;
        RECT 3.745 1.275 4.460 1.615 ;
        RECT 4.630 1.445 5.960 1.695 ;
        RECT 6.590 1.325 6.760 1.615 ;
        RECT 3.745 1.035 4.755 1.275 ;
        RECT 6.590 0.995 6.935 1.325 ;
        RECT 0.565 0.695 1.605 0.865 ;
        RECT 0.095 0.085 0.395 0.585 ;
        RECT 0.565 0.530 0.775 0.695 ;
        RECT 0.950 0.085 1.185 0.525 ;
        RECT 1.355 0.505 1.605 0.695 ;
        RECT 1.355 0.255 3.365 0.505 ;
        RECT 3.535 0.085 3.705 0.525 ;
        RECT 4.365 0.085 4.695 0.445 ;
        RECT 5.215 0.085 5.545 0.445 ;
        RECT 6.055 0.085 6.385 0.445 ;
        RECT 6.915 0.085 7.270 0.445 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 3.830 1.445 4.000 1.615 ;
        RECT 6.590 1.445 6.760 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
END sky130_fd_sc_hd__a211oi_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a221o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.970 1.075 2.300 1.275 ;
        RECT 1.970 0.675 2.255 1.075 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.470 1.075 2.835 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.225 1.075 1.700 1.275 ;
        RECT 1.420 0.675 1.700 1.075 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.610 1.075 1.055 1.275 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.440 1.285 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.660 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 3.320 1.795 3.575 2.465 ;
        RECT 3.405 0.665 3.575 1.795 ;
        RECT 3.390 0.585 3.575 0.665 ;
        RECT 3.320 0.255 3.575 0.585 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.175 1.625 0.345 2.465 ;
        RECT 0.515 2.295 1.685 2.465 ;
        RECT 0.515 1.795 0.845 2.295 ;
        RECT 1.355 2.255 1.685 2.295 ;
        RECT 1.875 2.215 2.230 2.635 ;
        RECT 1.015 2.035 1.245 2.125 ;
        RECT 2.400 2.035 2.650 2.465 ;
        RECT 1.015 1.795 2.650 2.035 ;
        RECT 2.820 1.875 3.150 2.635 ;
        RECT 0.175 1.455 3.235 1.625 ;
        RECT 3.065 0.905 3.235 1.455 ;
        RECT 0.175 0.735 1.240 0.905 ;
        RECT 0.175 0.255 0.345 0.735 ;
        RECT 0.515 0.085 0.845 0.565 ;
        RECT 1.070 0.505 1.240 0.735 ;
        RECT 2.435 0.735 3.235 0.905 ;
        RECT 2.435 0.505 2.605 0.735 ;
        RECT 1.070 0.255 2.605 0.505 ;
        RECT 2.775 0.085 3.105 0.565 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__a221o_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a221o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.970 1.075 2.300 1.275 ;
        RECT 1.970 0.675 2.255 1.075 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.470 1.075 2.835 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.225 1.075 1.700 1.275 ;
        RECT 1.420 0.675 1.700 1.075 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.610 1.075 1.055 1.275 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.440 1.285 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.105 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 3.320 1.795 3.575 2.465 ;
        RECT 3.405 0.665 3.575 1.795 ;
        RECT 3.390 0.585 3.575 0.665 ;
        RECT 3.320 0.255 3.575 0.585 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.175 1.625 0.345 2.465 ;
        RECT 0.515 2.295 1.685 2.465 ;
        RECT 0.515 1.795 0.845 2.295 ;
        RECT 1.355 2.255 1.685 2.295 ;
        RECT 1.875 2.215 2.230 2.635 ;
        RECT 1.015 2.035 1.245 2.125 ;
        RECT 2.400 2.035 2.650 2.465 ;
        RECT 1.015 1.795 2.650 2.035 ;
        RECT 2.820 1.875 3.150 2.635 ;
        RECT 0.175 1.455 3.235 1.625 ;
        RECT 3.065 0.905 3.235 1.455 ;
        RECT 3.745 1.445 3.915 2.635 ;
        RECT 0.175 0.735 1.240 0.905 ;
        RECT 0.175 0.255 0.345 0.735 ;
        RECT 0.515 0.085 0.845 0.565 ;
        RECT 1.070 0.505 1.240 0.735 ;
        RECT 2.435 0.735 3.235 0.905 ;
        RECT 2.435 0.505 2.605 0.735 ;
        RECT 1.070 0.255 2.605 0.505 ;
        RECT 2.775 0.085 3.105 0.565 ;
        RECT 3.745 0.085 3.915 0.980 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__a221o_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a221o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.855 1.105 4.060 1.285 ;
        RECT 2.855 1.075 3.190 1.105 ;
        RECT 3.710 1.075 4.060 1.105 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.265 1.075 2.680 1.285 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 5.235 1.075 6.035 1.285 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 6.270 1.075 7.280 1.285 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.230 1.075 4.725 1.285 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.435 1.015 ;
        RECT 0.155 -0.085 0.325 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.555 1.625 0.805 2.465 ;
        RECT 1.395 1.625 1.645 2.465 ;
        RECT 0.095 1.455 1.645 1.625 ;
        RECT 0.095 0.905 0.325 1.455 ;
        RECT 0.095 0.735 1.685 0.905 ;
        RECT 0.515 0.725 1.685 0.735 ;
        RECT 0.515 0.255 0.845 0.725 ;
        RECT 1.355 0.255 1.685 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.155 1.795 0.385 2.635 ;
        RECT 0.975 1.795 1.225 2.635 ;
        RECT 1.815 1.795 2.065 2.635 ;
        RECT 2.235 1.965 2.485 2.465 ;
        RECT 2.655 2.135 2.905 2.635 ;
        RECT 3.075 1.965 3.330 2.465 ;
        RECT 3.500 2.135 3.750 2.635 ;
        RECT 3.940 2.295 7.225 2.465 ;
        RECT 3.940 2.215 6.385 2.295 ;
        RECT 4.060 1.965 5.575 2.045 ;
        RECT 2.235 1.875 5.575 1.965 ;
        RECT 2.235 1.795 4.230 1.875 ;
        RECT 4.405 1.625 4.735 1.705 ;
        RECT 5.245 1.625 5.575 1.875 ;
        RECT 5.745 1.795 6.385 2.215 ;
        RECT 6.555 1.625 6.805 2.125 ;
        RECT 6.975 1.785 7.225 2.295 ;
        RECT 1.815 1.455 5.065 1.625 ;
        RECT 5.245 1.455 6.805 1.625 ;
        RECT 1.815 1.285 1.985 1.455 ;
        RECT 0.495 1.115 1.985 1.285 ;
        RECT 0.495 1.075 1.845 1.115 ;
        RECT 1.945 0.905 2.165 0.935 ;
        RECT 3.315 0.905 3.610 0.935 ;
        RECT 4.895 0.905 5.065 1.455 ;
        RECT 1.855 0.735 2.525 0.905 ;
        RECT 0.175 0.085 0.345 0.555 ;
        RECT 1.015 0.085 1.185 0.555 ;
        RECT 1.855 0.085 2.025 0.555 ;
        RECT 2.195 0.255 2.525 0.735 ;
        RECT 2.695 0.085 2.865 0.895 ;
        RECT 3.190 0.735 3.885 0.905 ;
        RECT 3.550 0.645 3.885 0.735 ;
        RECT 4.055 0.725 5.065 0.905 ;
        RECT 4.055 0.475 4.305 0.725 ;
        RECT 3.080 0.305 4.305 0.475 ;
        RECT 4.475 0.085 4.645 0.555 ;
        RECT 4.815 0.475 5.065 0.725 ;
        RECT 5.235 0.725 7.345 0.905 ;
        RECT 5.235 0.645 6.505 0.725 ;
        RECT 4.815 0.255 5.985 0.475 ;
        RECT 6.675 0.085 6.845 0.555 ;
        RECT 7.015 0.255 7.345 0.725 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 1.995 0.765 2.165 0.935 ;
        RECT 3.400 0.765 3.570 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
      LAYER met1 ;
        RECT 1.935 0.920 2.225 0.965 ;
        RECT 3.340 0.920 3.630 0.965 ;
        RECT 1.935 0.780 3.630 0.920 ;
        RECT 1.935 0.735 2.225 0.780 ;
        RECT 3.340 0.735 3.630 0.780 ;
  END
END sky130_fd_sc_hd__a221o_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a221oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.945 1.075 2.275 1.285 ;
        RECT 1.945 0.675 2.200 1.075 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.470 0.995 2.755 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.225 1.075 1.695 1.285 ;
        RECT 1.415 0.675 1.695 1.075 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.615 1.075 1.055 1.285 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.435 1.285 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.215 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.767000 ;
    PORT
      LAYER li1 ;
        RECT 0.175 1.625 0.345 2.465 ;
        RECT 2.150 1.625 3.135 1.665 ;
        RECT 0.175 1.495 3.135 1.625 ;
        RECT 0.175 1.455 2.300 1.495 ;
        RECT 0.170 0.735 1.235 0.905 ;
        RECT 2.925 0.825 3.135 1.495 ;
        RECT 0.170 0.255 0.345 0.735 ;
        RECT 1.065 0.505 1.235 0.735 ;
        RECT 2.380 0.655 3.135 0.825 ;
        RECT 2.380 0.505 2.580 0.655 ;
        RECT 1.065 0.255 2.580 0.505 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.515 2.295 1.685 2.465 ;
        RECT 0.515 1.795 0.765 2.295 ;
        RECT 1.355 2.255 1.685 2.295 ;
        RECT 1.875 2.215 2.205 2.635 ;
        RECT 1.015 2.045 1.240 2.125 ;
        RECT 2.375 2.045 2.625 2.465 ;
        RECT 1.015 1.835 2.625 2.045 ;
        RECT 2.795 1.875 3.125 2.635 ;
        RECT 1.015 1.795 2.025 1.835 ;
        RECT 0.515 0.085 0.845 0.565 ;
        RECT 2.750 0.085 3.080 0.485 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__a221oi_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a221oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.985 1.075 4.480 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.435 1.445 4.820 1.615 ;
        RECT 3.435 1.075 3.765 1.445 ;
        RECT 4.650 1.275 4.820 1.445 ;
        RECT 4.650 1.075 5.435 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.210 1.075 2.765 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.445 3.265 1.615 ;
        RECT 1.505 1.075 2.040 1.445 ;
        RECT 2.935 1.075 3.265 1.445 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.420 1.615 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.325 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.796500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.905 0.855 2.125 ;
        RECT 0.605 0.865 4.395 0.905 ;
        RECT 0.525 0.725 4.395 0.865 ;
        RECT 0.525 0.305 0.855 0.725 ;
        RECT 2.285 0.645 2.635 0.725 ;
        RECT 4.065 0.645 4.395 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.090 2.295 1.275 2.465 ;
        RECT 0.090 1.795 0.435 2.295 ;
        RECT 1.025 1.955 1.275 2.295 ;
        RECT 1.505 2.295 3.475 2.465 ;
        RECT 1.505 2.125 1.755 2.295 ;
        RECT 2.345 2.125 2.595 2.295 ;
        RECT 1.925 1.955 2.175 2.125 ;
        RECT 2.765 1.955 3.015 2.125 ;
        RECT 1.025 1.785 3.015 1.955 ;
        RECT 3.225 1.955 3.475 2.295 ;
        RECT 3.685 2.125 3.935 2.635 ;
        RECT 4.105 1.955 4.355 2.465 ;
        RECT 4.525 2.125 4.775 2.635 ;
        RECT 4.990 1.955 5.195 2.465 ;
        RECT 3.225 1.785 5.195 1.955 ;
        RECT 1.025 1.495 1.275 1.785 ;
        RECT 4.990 1.455 5.195 1.785 ;
        RECT 0.105 0.085 0.355 0.895 ;
        RECT 1.025 0.085 1.715 0.555 ;
        RECT 1.885 0.255 3.055 0.475 ;
        RECT 3.270 0.085 3.440 0.555 ;
        RECT 4.565 0.475 4.815 0.905 ;
        RECT 3.645 0.255 4.815 0.475 ;
        RECT 4.985 0.085 5.155 0.905 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__a221oi_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a221oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a221oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.475 1.075 7.885 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 5.965 1.445 8.265 1.615 ;
        RECT 5.965 1.075 6.295 1.445 ;
        RECT 8.095 1.275 8.265 1.445 ;
        RECT 8.095 1.075 9.575 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.935 0.995 5.285 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.595 1.445 5.795 1.615 ;
        RECT 3.595 1.325 3.765 1.445 ;
        RECT 3.415 0.995 3.765 1.325 ;
        RECT 5.465 1.075 5.795 1.445 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 1.335 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.535 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.593000 ;
    PORT
      LAYER li1 ;
        RECT 0.575 1.615 0.825 2.125 ;
        RECT 1.415 1.615 1.665 2.125 ;
        RECT 0.575 1.445 1.705 1.615 ;
        RECT 1.505 1.275 1.705 1.445 ;
        RECT 1.505 1.095 3.245 1.275 ;
        RECT 1.505 0.905 1.705 1.095 ;
        RECT 0.535 0.725 1.705 0.905 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 3.075 0.820 3.245 1.095 ;
        RECT 5.510 0.820 6.460 0.905 ;
        RECT 3.075 0.735 7.765 0.820 ;
        RECT 3.075 0.645 5.680 0.735 ;
        RECT 6.290 0.645 7.765 0.735 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.090 2.295 2.125 2.465 ;
        RECT 0.090 1.445 0.405 2.295 ;
        RECT 0.995 1.785 1.245 2.295 ;
        RECT 1.875 1.615 2.125 2.295 ;
        RECT 2.315 2.215 6.005 2.465 ;
        RECT 6.175 2.215 8.185 2.635 ;
        RECT 2.315 1.795 2.565 2.215 ;
        RECT 5.755 2.045 6.005 2.215 ;
        RECT 8.355 2.045 8.525 2.465 ;
        RECT 2.735 1.835 5.585 2.045 ;
        RECT 2.735 1.615 3.030 1.835 ;
        RECT 5.755 1.785 8.605 2.045 ;
        RECT 8.775 1.795 8.945 2.635 ;
        RECT 1.875 1.445 3.030 1.615 ;
        RECT 8.435 1.615 8.605 1.785 ;
        RECT 9.155 1.615 9.405 2.465 ;
        RECT 8.435 1.445 9.405 1.615 ;
        RECT 0.115 0.085 0.365 0.895 ;
        RECT 1.875 0.645 2.905 0.925 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.645 ;
        RECT 2.735 0.595 2.905 0.645 ;
        RECT 7.935 0.725 9.025 0.905 ;
        RECT 2.235 0.425 2.610 0.475 ;
        RECT 3.035 0.425 5.585 0.475 ;
        RECT 2.235 0.255 5.585 0.425 ;
        RECT 5.835 0.085 6.005 0.555 ;
        RECT 7.935 0.475 8.185 0.725 ;
        RECT 6.175 0.255 8.185 0.475 ;
        RECT 8.355 0.085 8.525 0.555 ;
        RECT 8.695 0.255 9.025 0.725 ;
        RECT 9.195 0.085 9.365 0.905 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
  END
END sky130_fd_sc_hd__a221oi_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a222oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a222oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.615 1.000 2.925 1.330 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 3.095 1.000 3.435 1.330 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 2.135 1.000 2.445 1.330 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 1.655 1.000 1.965 1.330 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.000 0.545 1.315 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 0.715 1.000 1.085 1.315 ;
    END
  END C2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.240 3.675 1.005 ;
        RECT 0.000 0.000 3.680 0.240 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER li1 ;
        RECT 0.095 2.255 0.425 2.465 ;
        RECT 0.095 1.680 0.345 2.255 ;
        RECT 0.095 1.670 0.425 1.680 ;
        RECT 1.015 1.670 1.185 1.830 ;
        RECT 0.095 1.500 1.425 1.670 ;
        RECT 0.095 1.485 0.425 1.500 ;
        RECT 1.255 1.330 1.425 1.500 ;
        RECT 1.255 0.815 1.480 1.330 ;
        RECT 0.095 0.645 2.645 0.815 ;
        RECT 0.095 0.255 0.425 0.645 ;
        RECT 2.315 0.295 2.645 0.645 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.595 2.295 2.185 2.465 ;
        RECT 0.595 2.075 0.765 2.295 ;
        RECT 2.015 2.135 2.185 2.295 ;
        RECT 2.355 2.255 2.685 2.465 ;
        RECT 0.515 1.875 0.845 2.075 ;
        RECT 1.515 1.980 1.915 1.995 ;
        RECT 1.515 1.970 1.935 1.980 ;
        RECT 1.515 1.965 1.970 1.970 ;
        RECT 1.515 1.825 2.015 1.965 ;
        RECT 2.355 1.825 2.605 2.255 ;
        RECT 2.855 2.075 3.025 2.635 ;
        RECT 3.255 2.255 3.595 2.465 ;
        RECT 2.775 1.905 3.105 2.075 ;
        RECT 1.845 1.735 2.605 1.825 ;
        RECT 3.335 1.735 3.595 2.255 ;
        RECT 1.845 1.670 2.685 1.735 ;
        RECT 3.220 1.670 3.595 1.735 ;
        RECT 1.845 1.655 3.595 1.670 ;
        RECT 2.355 1.500 3.595 1.655 ;
        RECT 0.875 0.085 1.605 0.465 ;
        RECT 3.255 0.085 3.585 0.815 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__a222oi_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a311o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.965 0.995 2.310 1.325 ;
        RECT 1.965 0.765 2.155 0.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.510 0.750 1.705 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.905 0.995 1.240 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.620 0.995 3.095 1.325 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.350 0.995 3.535 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.675 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.454000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.785 0.425 2.425 ;
        RECT 0.085 0.670 0.255 1.785 ;
        RECT 0.085 0.255 0.395 0.670 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.595 2.175 0.840 2.635 ;
        RECT 1.015 2.005 1.265 2.465 ;
        RECT 1.455 2.255 2.125 2.635 ;
        RECT 2.325 2.005 2.575 2.465 ;
        RECT 1.015 1.835 2.575 2.005 ;
        RECT 3.335 1.665 3.505 2.465 ;
        RECT 0.565 1.495 3.505 1.665 ;
        RECT 0.565 1.325 0.735 1.495 ;
        RECT 0.425 0.995 0.735 1.325 ;
        RECT 0.565 0.825 0.735 0.995 ;
        RECT 0.565 0.655 1.260 0.825 ;
        RECT 0.590 0.085 0.920 0.465 ;
        RECT 1.090 0.425 1.260 0.655 ;
        RECT 2.325 0.655 3.505 0.825 ;
        RECT 2.325 0.425 2.495 0.655 ;
        RECT 1.090 0.255 2.495 0.425 ;
        RECT 2.765 0.085 3.095 0.485 ;
        RECT 3.335 0.255 3.505 0.655 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__a311o_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a311o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.440 0.995 2.675 1.325 ;
        RECT 2.440 0.605 2.620 0.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.895 0.605 2.165 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.495 0.995 1.710 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.895 0.995 3.235 1.325 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.695 0.995 4.005 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.135 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.295 0.845 2.425 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.160 1.835 1.380 2.635 ;
        RECT 1.590 2.005 1.840 2.465 ;
        RECT 2.125 2.255 2.455 2.635 ;
        RECT 2.715 2.005 3.025 2.465 ;
        RECT 1.590 1.835 3.025 2.005 ;
        RECT 3.795 1.665 3.965 2.465 ;
        RECT 1.015 1.495 3.965 1.665 ;
        RECT 0.090 0.085 0.345 0.885 ;
        RECT 1.015 0.825 1.185 1.495 ;
        RECT 1.015 0.655 1.695 0.825 ;
        RECT 1.015 0.085 1.345 0.465 ;
        RECT 1.525 0.425 1.695 0.655 ;
        RECT 2.790 0.655 3.965 0.825 ;
        RECT 2.790 0.425 2.960 0.655 ;
        RECT 1.525 0.255 2.960 0.425 ;
        RECT 3.220 0.085 3.550 0.485 ;
        RECT 3.795 0.255 3.965 0.655 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__a311o_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a311o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 6.945 1.075 7.275 1.615 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 5.255 1.075 6.040 1.285 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.515 1.075 4.945 1.285 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.060 1.285 1.255 1.625 ;
        RECT 1.060 1.075 1.505 1.285 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.745 0.350 1.625 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.355 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.904000 ;
    PORT
      LAYER li1 ;
        RECT 2.715 1.545 3.885 1.715 ;
        RECT 2.910 0.885 3.105 1.545 ;
        RECT 2.295 0.715 3.305 0.885 ;
        RECT 2.295 0.465 2.465 0.715 ;
        RECT 3.135 0.465 3.305 0.715 ;
        RECT 2.195 0.295 2.545 0.465 ;
        RECT 3.055 0.295 3.385 0.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.175 2.295 2.025 2.465 ;
        RECT 0.175 1.795 0.345 2.295 ;
        RECT 0.515 1.955 0.845 2.125 ;
        RECT 0.595 0.885 0.765 1.955 ;
        RECT 1.015 1.795 1.185 2.295 ;
        RECT 1.435 1.625 1.605 2.125 ;
        RECT 1.855 1.795 2.025 2.295 ;
        RECT 2.295 2.255 2.625 2.635 ;
        RECT 3.135 2.255 3.465 2.635 ;
        RECT 3.975 2.255 4.305 2.635 ;
        RECT 4.475 2.085 4.645 2.465 ;
        RECT 4.815 2.255 5.175 2.635 ;
        RECT 5.375 2.085 5.545 2.465 ;
        RECT 5.715 2.255 6.045 2.635 ;
        RECT 6.595 2.085 6.765 2.465 ;
        RECT 2.195 1.915 6.765 2.085 ;
        RECT 2.195 1.625 2.385 1.915 ;
        RECT 4.475 1.795 4.645 1.915 ;
        RECT 5.375 1.795 5.545 1.915 ;
        RECT 6.595 1.795 6.765 1.915 ;
        RECT 6.935 1.795 7.270 2.635 ;
        RECT 1.435 1.455 2.385 1.625 ;
        RECT 4.150 1.455 6.685 1.625 ;
        RECT 4.150 1.245 4.320 1.455 ;
        RECT 1.855 1.075 2.705 1.245 ;
        RECT 3.275 1.075 4.320 1.245 ;
        RECT 1.855 0.885 2.025 1.075 ;
        RECT 0.595 0.715 2.025 0.885 ;
        RECT 4.355 0.715 6.005 0.885 ;
        RECT 0.095 0.085 0.345 0.565 ;
        RECT 0.595 0.465 0.765 0.715 ;
        RECT 0.515 0.295 0.845 0.465 ;
        RECT 1.015 0.085 1.185 0.545 ;
        RECT 1.435 0.465 1.605 0.715 ;
        RECT 1.355 0.295 1.685 0.465 ;
        RECT 1.855 0.085 2.025 0.545 ;
        RECT 2.715 0.085 2.885 0.545 ;
        RECT 3.555 0.085 4.065 0.545 ;
        RECT 4.355 0.465 4.525 0.715 ;
        RECT 5.675 0.645 6.005 0.715 ;
        RECT 4.275 0.295 4.605 0.465 ;
        RECT 4.775 0.085 4.945 0.545 ;
        RECT 6.175 0.465 6.345 0.885 ;
        RECT 6.515 0.825 6.685 1.455 ;
        RECT 6.515 0.645 6.845 0.825 ;
        RECT 7.015 0.500 7.270 0.905 ;
        RECT 5.255 0.425 6.345 0.465 ;
        RECT 6.935 0.425 7.270 0.500 ;
        RECT 5.255 0.255 7.270 0.425 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
END sky130_fd_sc_hd__a311o_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a311oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.195 0.995 1.455 1.325 ;
        RECT 1.195 0.660 1.365 0.995 ;
        RECT 0.965 0.265 1.365 0.660 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.600 0.995 1.025 1.325 ;
        RECT 0.600 0.265 0.795 0.995 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.420 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.950 2.005 2.230 2.355 ;
        RECT 1.710 1.835 2.230 2.005 ;
        RECT 1.710 0.995 1.935 1.835 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.995 2.685 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.790 1.015 ;
        RECT 0.155 -0.085 0.325 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.659750 ;
    PORT
      LAYER li1 ;
        RECT 2.410 1.665 2.650 2.335 ;
        RECT 2.105 1.495 2.650 1.665 ;
        RECT 2.105 0.825 2.275 1.495 ;
        RECT 1.535 0.655 2.650 0.825 ;
        RECT 1.535 0.255 1.705 0.655 ;
        RECT 2.405 0.295 2.650 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.095 1.495 0.425 2.635 ;
        RECT 0.600 1.745 0.770 2.305 ;
        RECT 0.940 1.915 1.200 2.635 ;
        RECT 1.370 2.175 1.700 2.345 ;
        RECT 1.370 1.745 1.540 2.175 ;
        RECT 0.600 1.575 1.540 1.745 ;
        RECT 0.095 0.085 0.425 0.805 ;
        RECT 1.905 0.085 2.235 0.485 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__a311oi_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a311oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.000 0.995 3.115 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.055 0.995 1.805 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.995 0.800 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.395 0.995 4.055 1.325 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 5.175 1.295 5.410 1.625 ;
        RECT 4.730 1.075 5.410 1.295 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.515 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.141000 ;
    PORT
      LAYER li1 ;
        RECT 4.660 1.915 5.005 2.085 ;
        RECT 4.660 1.745 4.990 1.915 ;
        RECT 4.660 1.680 5.005 1.745 ;
        RECT 4.260 1.575 5.005 1.680 ;
        RECT 4.260 1.510 4.990 1.575 ;
        RECT 4.260 0.825 4.475 1.510 ;
        RECT 2.295 0.655 5.345 0.825 ;
        RECT 3.235 0.255 3.405 0.655 ;
        RECT 4.085 0.255 4.255 0.655 ;
        RECT 5.175 0.255 5.345 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.095 1.495 0.345 2.635 ;
        RECT 0.595 1.745 0.765 2.465 ;
        RECT 0.935 1.915 1.265 2.635 ;
        RECT 1.435 1.745 1.605 2.465 ;
        RECT 1.785 1.915 2.135 2.635 ;
        RECT 2.305 1.745 2.475 2.465 ;
        RECT 2.645 1.915 2.975 2.635 ;
        RECT 4.110 2.425 4.440 2.465 ;
        RECT 5.175 2.425 5.345 2.465 ;
        RECT 3.145 2.255 5.345 2.425 ;
        RECT 3.585 1.745 3.915 2.085 ;
        RECT 4.110 1.915 4.440 2.255 ;
        RECT 5.175 1.795 5.345 2.255 ;
        RECT 0.595 1.575 3.915 1.745 ;
        RECT 0.175 0.655 2.105 0.825 ;
        RECT 0.175 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.255 1.185 0.655 ;
        RECT 1.355 0.305 3.045 0.475 ;
        RECT 3.585 0.085 3.915 0.465 ;
        RECT 4.675 0.085 5.005 0.465 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__a311oi_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a311oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a311oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.805 0.995 5.420 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.935 0.995 3.550 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.120 0.995 1.735 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 5.670 0.995 6.855 1.630 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 7.935 0.995 9.530 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.655 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.898500 ;
    PORT
      LAYER li1 ;
        RECT 7.415 1.715 7.735 1.975 ;
        RECT 7.975 1.715 8.305 2.085 ;
        RECT 8.815 1.715 9.145 2.085 ;
        RECT 7.415 1.545 9.145 1.715 ;
        RECT 7.415 0.805 7.735 1.545 ;
        RECT 7.975 1.530 8.305 1.545 ;
        RECT 3.975 0.635 9.485 0.805 ;
        RECT 6.575 0.255 6.745 0.635 ;
        RECT 7.415 0.255 7.585 0.635 ;
        RECT 8.475 0.255 8.645 0.635 ;
        RECT 9.315 0.255 9.485 0.635 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.095 1.575 0.425 2.635 ;
        RECT 0.595 1.665 0.765 2.465 ;
        RECT 0.935 1.915 1.265 2.635 ;
        RECT 1.435 1.665 1.605 2.465 ;
        RECT 1.775 1.915 2.105 2.635 ;
        RECT 2.275 1.665 2.445 2.465 ;
        RECT 2.615 1.915 2.945 2.635 ;
        RECT 3.115 1.665 3.285 2.465 ;
        RECT 3.455 1.915 3.785 2.635 ;
        RECT 3.955 1.665 4.125 2.465 ;
        RECT 4.295 1.915 4.625 2.635 ;
        RECT 4.795 2.085 4.965 2.465 ;
        RECT 5.135 2.255 5.465 2.635 ;
        RECT 5.655 2.255 9.565 2.425 ;
        RECT 4.795 1.915 7.245 2.085 ;
        RECT 4.795 1.665 4.965 1.915 ;
        RECT 9.315 1.835 9.565 2.255 ;
        RECT 0.595 1.495 4.965 1.665 ;
        RECT 0.175 0.635 3.785 0.805 ;
        RECT 0.175 0.255 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.255 1.185 0.635 ;
        RECT 1.355 0.085 1.685 0.465 ;
        RECT 1.855 0.255 2.025 0.635 ;
        RECT 2.195 0.295 5.565 0.465 ;
        RECT 6.075 0.085 6.405 0.465 ;
        RECT 6.915 0.085 7.245 0.465 ;
        RECT 7.975 0.085 8.305 0.465 ;
        RECT 8.815 0.085 9.145 0.465 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
  END
END sky130_fd_sc_hd__a311oi_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a2111o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111o_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.995 3.290 1.325 ;
        RECT 2.985 0.845 3.290 0.995 ;
        RECT 2.985 0.285 3.540 0.845 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.510 1.025 4.010 1.290 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.400 0.995 2.680 2.465 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.890 1.050 2.220 2.465 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.290 1.720 2.465 ;
        RECT 1.290 1.050 1.720 1.290 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.125 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
        RECT 1.985 -0.085 2.155 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504500 ;
    PORT
      LAYER li1 ;
        RECT 0.135 1.620 0.390 2.460 ;
        RECT 0.135 0.255 0.465 1.620 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.565 1.815 0.895 2.635 ;
        RECT 1.135 1.645 1.345 2.460 ;
        RECT 0.695 1.465 1.345 1.645 ;
        RECT 2.860 1.665 3.145 2.460 ;
        RECT 3.325 1.835 3.540 2.635 ;
        RECT 3.720 1.665 3.990 2.460 ;
        RECT 2.860 1.495 3.990 1.665 ;
        RECT 0.695 0.825 0.915 1.465 ;
        RECT 0.695 0.655 2.805 0.825 ;
        RECT 0.695 0.650 1.915 0.655 ;
        RECT 0.635 0.085 1.310 0.470 ;
        RECT 1.585 0.260 1.915 0.650 ;
        RECT 2.085 0.085 2.430 0.485 ;
        RECT 2.600 0.260 2.805 0.655 ;
        RECT 3.715 0.085 3.955 0.760 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__a2111o_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a2111o_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111o_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.365 0.955 3.775 1.740 ;
        RECT 3.505 0.825 3.775 0.955 ;
        RECT 3.505 0.290 3.995 0.825 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.945 0.995 4.515 1.740 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.905 0.995 3.195 1.740 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.425 0.995 2.735 2.355 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.960 1.325 2.255 2.355 ;
        RECT 1.885 0.995 2.255 1.325 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.095 0.105 4.585 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.255 0.895 2.390 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.085 1.635 0.435 2.635 ;
        RECT 1.065 1.495 1.315 2.635 ;
        RECT 1.495 1.495 1.785 2.465 ;
        RECT 3.070 2.085 3.400 2.465 ;
        RECT 3.590 2.255 3.920 2.635 ;
        RECT 4.090 2.085 4.515 2.465 ;
        RECT 3.070 1.915 4.515 2.085 ;
        RECT 1.495 1.325 1.705 1.495 ;
        RECT 1.065 1.075 1.705 1.325 ;
        RECT 0.085 0.085 0.435 0.885 ;
        RECT 1.065 0.445 1.325 0.865 ;
        RECT 1.495 0.785 1.705 1.075 ;
        RECT 1.495 0.615 3.335 0.785 ;
        RECT 1.065 0.085 2.010 0.445 ;
        RECT 2.180 0.255 2.420 0.615 ;
        RECT 2.590 0.085 2.920 0.445 ;
        RECT 3.090 0.255 3.335 0.615 ;
        RECT 4.165 0.085 4.515 0.805 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__a2111o_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a2111o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111o_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.825 1.075 4.495 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.675 1.075 5.625 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.450 0.975 3.255 1.285 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.040 0.975 2.280 1.285 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.370 1.625 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.090 0.105 7.805 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER li1 ;
        RECT 6.165 1.715 6.355 2.465 ;
        RECT 7.025 1.715 7.215 2.465 ;
        RECT 6.165 1.635 7.215 1.715 ;
        RECT 6.165 1.465 7.735 1.635 ;
        RECT 7.490 0.805 7.735 1.465 ;
        RECT 6.165 0.635 7.735 0.805 ;
        RECT 6.165 0.255 6.355 0.635 ;
        RECT 7.025 0.255 7.215 0.635 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.110 2.295 2.160 2.465 ;
        RECT 0.110 1.795 0.370 2.295 ;
        RECT 0.540 0.805 0.870 2.125 ;
        RECT 1.040 1.455 1.230 2.295 ;
        RECT 1.400 1.625 1.730 2.125 ;
        RECT 1.900 1.795 2.160 2.295 ;
        RECT 2.340 2.295 3.650 2.465 ;
        RECT 2.340 1.795 2.675 2.295 ;
        RECT 2.845 1.625 3.100 2.125 ;
        RECT 3.320 1.995 3.650 2.295 ;
        RECT 3.865 2.165 4.195 2.635 ;
        RECT 4.365 1.995 4.625 2.415 ;
        RECT 4.805 2.255 5.140 2.635 ;
        RECT 5.310 1.995 5.495 2.465 ;
        RECT 3.320 1.795 5.495 1.995 ;
        RECT 5.665 1.800 5.995 2.635 ;
        RECT 6.525 1.885 6.855 2.635 ;
        RECT 7.385 1.805 7.715 2.635 ;
        RECT 1.400 1.455 3.100 1.625 ;
        RECT 3.465 1.445 5.975 1.625 ;
        RECT 3.465 0.805 3.655 1.445 ;
        RECT 5.795 1.245 5.975 1.445 ;
        RECT 5.795 1.075 7.320 1.245 ;
        RECT 0.180 0.635 3.655 0.805 ;
        RECT 0.180 0.255 0.440 0.635 ;
        RECT 1.110 0.615 3.655 0.635 ;
        RECT 3.825 0.615 5.495 0.785 ;
        RECT 0.610 0.085 0.940 0.465 ;
        RECT 1.110 0.255 1.340 0.615 ;
        RECT 1.510 0.085 1.840 0.445 ;
        RECT 2.015 0.255 2.240 0.615 ;
        RECT 3.465 0.445 3.655 0.615 ;
        RECT 2.420 0.085 3.295 0.445 ;
        RECT 3.465 0.255 4.585 0.445 ;
        RECT 4.805 0.085 5.140 0.445 ;
        RECT 5.310 0.255 5.495 0.615 ;
        RECT 5.665 0.085 5.995 0.515 ;
        RECT 6.525 0.085 6.855 0.445 ;
        RECT 7.385 0.085 7.715 0.465 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
  END
END sky130_fd_sc_hd__a2111o_4

#--------EOF---------

MACRO sky130_fd_sc_hd__a2111oi_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.355 1.400 2.625 1.735 ;
        RECT 2.035 1.070 2.625 1.400 ;
        RECT 2.355 0.660 2.625 1.070 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.795 0.650 3.135 1.735 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.495 1.055 1.845 1.735 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.055 1.325 2.360 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.730 0.435 1.655 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.195 0.105 2.910 0.785 ;
        RECT 0.195 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.424000 ;
    PORT
      LAYER li1 ;
        RECT 0.360 1.825 0.785 2.465 ;
        RECT 0.605 0.885 0.785 1.825 ;
        RECT 0.605 0.635 2.040 0.885 ;
        RECT 0.785 0.615 2.040 0.635 ;
        RECT 0.785 0.255 1.040 0.615 ;
        RECT 1.710 0.280 2.040 0.615 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 1.540 2.085 1.870 2.465 ;
        RECT 2.040 2.255 2.370 2.635 ;
        RECT 2.540 2.085 2.870 2.465 ;
        RECT 1.540 1.905 2.870 2.085 ;
        RECT 0.285 0.085 0.615 0.465 ;
        RECT 1.210 0.085 1.540 0.445 ;
        RECT 2.470 0.085 2.800 0.480 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__a2111oi_0

#--------EOF---------

MACRO sky130_fd_sc_hd__a2111oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.440 0.995 2.725 1.400 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.020 3.540 1.290 ;
        RECT 2.905 0.350 3.090 1.020 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.940 1.400 2.215 2.455 ;
        RECT 1.940 1.050 2.270 1.400 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.435 1.050 1.770 2.455 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.785 1.050 1.235 2.455 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.105 3.675 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
        RECT 1.975 -0.065 2.145 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.388750 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.880 0.530 2.460 ;
        RECT 0.145 0.815 2.300 0.880 ;
        RECT 0.145 0.705 2.420 0.815 ;
        RECT 0.145 0.700 1.375 0.705 ;
        RECT 1.045 0.260 1.375 0.700 ;
        RECT 2.090 0.305 2.420 0.705 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 2.395 1.750 2.625 2.460 ;
        RECT 2.800 1.920 3.130 2.635 ;
        RECT 3.310 1.750 3.505 2.460 ;
        RECT 2.395 1.580 3.505 1.750 ;
        RECT 0.315 0.085 0.630 0.525 ;
        RECT 1.550 0.085 1.880 0.535 ;
        RECT 3.270 0.085 3.510 0.760 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__a2111oi_1

#--------EOF---------

MACRO sky130_fd_sc_hd__a2111oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.465 1.445 5.290 1.675 ;
        RECT 3.465 0.985 3.715 1.445 ;
        RECT 4.895 0.995 5.290 1.445 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.970 1.015 4.725 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.185 1.030 2.855 1.275 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 1.445 1.800 1.680 ;
        RECT 0.125 1.045 0.455 1.445 ;
        RECT 1.615 1.275 1.800 1.445 ;
        RECT 1.615 1.030 1.975 1.275 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.755 1.075 1.425 1.275 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.105 5.440 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.212750 ;
    PORT
      LAYER li1 ;
        RECT 0.900 1.850 2.140 2.105 ;
        RECT 1.970 1.625 2.140 1.850 ;
        RECT 1.970 1.445 3.255 1.625 ;
        RECT 3.025 0.845 3.255 1.445 ;
        RECT 0.120 0.805 3.255 0.845 ;
        RECT 0.120 0.615 5.355 0.805 ;
        RECT 0.120 0.255 0.380 0.615 ;
        RECT 1.050 0.255 1.295 0.615 ;
        RECT 1.965 0.255 2.295 0.615 ;
        RECT 2.965 0.275 3.295 0.615 ;
        RECT 5.020 0.295 5.355 0.615 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.100 2.295 2.985 2.465 ;
        RECT 0.100 2.275 2.185 2.295 ;
        RECT 0.100 1.870 0.460 2.275 ;
        RECT 2.815 2.135 2.985 2.295 ;
        RECT 3.155 2.095 3.520 2.465 ;
        RECT 3.690 2.275 4.020 2.635 ;
        RECT 4.190 2.105 4.400 2.465 ;
        RECT 4.570 2.275 4.900 2.635 ;
        RECT 5.070 2.105 5.400 2.465 ;
        RECT 4.190 2.095 5.400 2.105 ;
        RECT 2.310 1.965 2.640 2.060 ;
        RECT 3.155 1.965 5.400 2.095 ;
        RECT 2.310 1.845 5.400 1.965 ;
        RECT 2.310 1.795 3.335 1.845 ;
        RECT 0.550 0.085 0.880 0.445 ;
        RECT 1.465 0.085 1.795 0.445 ;
        RECT 2.465 0.085 2.795 0.445 ;
        RECT 4.125 0.085 4.455 0.445 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__a2111oi_2

#--------EOF---------

MACRO sky130_fd_sc_hd__a2111oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__a2111oi_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.095 1.020 7.745 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 7.960 1.020 9.990 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.955 1.020 5.650 1.275 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 2.055 1.020 3.745 1.275 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.495 1.020 1.845 1.275 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.955 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.009500 ;
    PORT
      LAYER li1 ;
        RECT 0.530 1.685 0.860 2.085 ;
        RECT 1.390 1.685 1.720 2.085 ;
        RECT 0.530 1.655 1.720 1.685 ;
        RECT 0.145 1.475 1.720 1.655 ;
        RECT 0.145 0.785 0.320 1.475 ;
        RECT 0.145 0.615 7.620 0.785 ;
        RECT 0.615 0.455 0.790 0.615 ;
        RECT 1.460 0.455 1.650 0.615 ;
        RECT 2.400 0.455 2.590 0.615 ;
        RECT 3.260 0.455 3.510 0.615 ;
        RECT 4.180 0.455 4.420 0.615 ;
        RECT 5.090 0.455 5.275 0.615 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.100 2.255 3.870 2.445 ;
        RECT 0.100 1.835 0.360 2.255 ;
        RECT 1.030 1.855 1.220 2.255 ;
        RECT 1.890 1.855 2.080 2.255 ;
        RECT 2.250 1.685 2.580 2.085 ;
        RECT 2.750 1.855 2.940 2.255 ;
        RECT 3.110 1.685 3.440 2.085 ;
        RECT 3.610 1.835 3.870 2.255 ;
        RECT 4.060 2.275 6.050 2.445 ;
        RECT 4.060 2.255 5.180 2.275 ;
        RECT 4.060 1.835 4.320 2.255 ;
        RECT 2.250 1.655 3.440 1.685 ;
        RECT 4.490 1.685 4.820 2.085 ;
        RECT 4.990 1.855 5.180 2.255 ;
        RECT 5.350 1.685 5.680 2.085 ;
        RECT 4.490 1.655 5.680 1.685 ;
        RECT 2.250 1.475 5.680 1.655 ;
        RECT 5.860 1.615 6.050 2.275 ;
        RECT 6.220 1.785 6.550 2.635 ;
        RECT 6.720 1.615 6.910 2.315 ;
        RECT 7.080 1.805 7.410 2.635 ;
        RECT 7.580 1.665 7.910 2.315 ;
        RECT 8.080 1.895 8.410 2.635 ;
        RECT 8.580 1.670 8.840 2.290 ;
        RECT 9.030 1.915 9.360 2.635 ;
        RECT 9.530 1.670 9.770 2.260 ;
        RECT 8.580 1.665 9.770 1.670 ;
        RECT 7.580 1.615 9.770 1.665 ;
        RECT 5.860 1.445 9.770 1.615 ;
        RECT 7.885 0.615 9.865 0.785 ;
        RECT 7.885 0.445 8.075 0.615 ;
        RECT 0.115 0.085 0.445 0.445 ;
        RECT 0.960 0.085 1.290 0.445 ;
        RECT 1.820 0.085 2.230 0.445 ;
        RECT 2.760 0.085 3.090 0.445 ;
        RECT 3.680 0.085 4.010 0.445 ;
        RECT 4.590 0.085 4.920 0.445 ;
        RECT 5.445 0.085 5.780 0.445 ;
        RECT 5.980 0.275 8.075 0.445 ;
        RECT 8.245 0.085 8.575 0.445 ;
        RECT 8.745 0.300 8.935 0.615 ;
        RECT 9.105 0.085 9.435 0.445 ;
        RECT 9.605 0.290 9.865 0.615 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
  END
END sky130_fd_sc_hd__a2111oi_4

#--------EOF---------

MACRO sky130_fd_sc_hd__and2_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.185 0.430 1.955 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.940 1.080 1.270 1.615 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.070 0.105 1.980 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.280900 ;
    PORT
      LAYER li1 ;
        RECT 1.790 1.835 2.215 2.465 ;
        RECT 1.950 0.525 2.215 1.835 ;
        RECT 1.560 0.255 2.215 0.525 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.160 2.175 0.430 2.635 ;
        RECT 0.600 2.135 0.865 2.465 ;
        RECT 0.600 0.950 0.770 2.135 ;
        RECT 1.110 1.835 1.620 2.635 ;
        RECT 0.185 0.910 0.770 0.950 ;
        RECT 1.450 0.910 1.780 1.435 ;
        RECT 0.185 0.695 1.780 0.910 ;
        RECT 0.185 0.280 0.490 0.695 ;
        RECT 0.950 0.085 1.390 0.525 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__and2_0

#--------EOF---------

MACRO sky130_fd_sc_hd__and2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.325 0.365 1.685 ;
        RECT 0.100 1.075 0.775 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.075 1.335 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.145 0.925 2.095 1.015 ;
        RECT 0.165 0.105 2.095 0.925 ;
        RECT 0.165 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.657000 ;
    PORT
      LAYER li1 ;
        RECT 1.755 1.915 2.215 2.465 ;
        RECT 1.965 0.545 2.215 1.915 ;
        RECT 1.655 0.255 2.215 0.545 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.285 1.965 0.565 2.635 ;
        RECT 0.735 1.745 1.035 2.295 ;
        RECT 1.235 1.915 1.565 2.635 ;
        RECT 0.735 1.575 1.675 1.745 ;
        RECT 1.505 1.325 1.675 1.575 ;
        RECT 1.505 0.995 1.795 1.325 ;
        RECT 1.505 0.905 1.675 0.995 ;
        RECT 0.285 0.715 1.675 0.905 ;
        RECT 0.285 0.355 0.615 0.715 ;
        RECT 1.235 0.085 1.485 0.545 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__and2_1

#--------EOF---------

MACRO sky130_fd_sc_hd__and2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.325 0.400 1.765 ;
        RECT 0.085 1.075 0.775 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.075 1.335 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.155 0.925 2.745 1.015 ;
        RECT 0.175 0.105 2.745 0.925 ;
        RECT 0.175 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.643500 ;
    PORT
      LAYER li1 ;
        RECT 1.765 1.915 2.215 2.465 ;
        RECT 1.965 0.545 2.215 1.915 ;
        RECT 1.665 0.255 2.215 0.545 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.285 1.965 0.565 2.635 ;
        RECT 0.735 1.745 1.035 2.295 ;
        RECT 1.245 1.915 1.575 2.635 ;
        RECT 0.735 1.575 1.675 1.745 ;
        RECT 1.505 1.325 1.675 1.575 ;
        RECT 2.385 1.495 2.675 2.635 ;
        RECT 1.505 0.995 1.795 1.325 ;
        RECT 1.505 0.905 1.675 0.995 ;
        RECT 0.285 0.715 1.675 0.905 ;
        RECT 0.285 0.355 0.615 0.715 ;
        RECT 1.245 0.085 1.495 0.545 ;
        RECT 2.385 0.085 2.675 0.885 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__and2_2

#--------EOF---------

MACRO sky130_fd_sc_hd__and2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.995 0.435 1.615 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.995 0.980 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.190 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER li1 ;
        RECT 1.530 1.760 1.720 2.465 ;
        RECT 2.390 1.765 2.580 2.465 ;
        RECT 2.390 1.760 3.135 1.765 ;
        RECT 1.530 1.535 3.135 1.760 ;
        RECT 2.855 0.845 3.135 1.535 ;
        RECT 1.530 0.615 3.135 0.845 ;
        RECT 1.530 0.515 1.720 0.615 ;
        RECT 2.390 0.255 2.580 0.615 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.095 1.880 0.425 2.635 ;
        RECT 0.605 1.750 0.785 2.465 ;
        RECT 0.990 1.935 1.320 2.635 ;
        RECT 1.890 1.935 2.220 2.635 ;
        RECT 2.750 1.935 3.080 2.635 ;
        RECT 0.605 1.580 1.360 1.750 ;
        RECT 1.150 1.355 1.360 1.580 ;
        RECT 1.150 1.020 2.685 1.355 ;
        RECT 1.150 0.805 1.360 1.020 ;
        RECT 0.095 0.615 1.360 0.805 ;
        RECT 0.095 0.255 0.425 0.615 ;
        RECT 0.955 0.085 1.285 0.445 ;
        RECT 1.890 0.085 2.220 0.445 ;
        RECT 2.750 0.085 3.080 0.445 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__and2_4

#--------EOF---------

MACRO sky130_fd_sc_hd__and2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.445 1.615 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.480 1.645 2.175 1.955 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.825 0.785 2.755 1.015 ;
        RECT 0.005 0.105 2.755 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 2.350 1.580 2.655 2.365 ;
        RECT 2.480 0.775 2.655 1.580 ;
        RECT 2.415 0.255 2.655 0.775 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.175 2.015 0.345 2.445 ;
        RECT 0.515 2.185 0.845 2.635 ;
        RECT 0.175 1.785 0.850 2.015 ;
        RECT 0.615 1.135 0.850 1.785 ;
        RECT 1.020 1.475 1.305 2.420 ;
        RECT 1.485 2.165 2.170 2.635 ;
        RECT 1.020 1.325 1.880 1.475 ;
        RECT 1.020 1.305 2.305 1.325 ;
        RECT 0.615 0.805 1.150 1.135 ;
        RECT 1.320 0.945 2.305 1.305 ;
        RECT 0.615 0.655 0.835 0.805 ;
        RECT 0.090 0.085 0.425 0.590 ;
        RECT 0.595 0.280 0.835 0.655 ;
        RECT 1.320 0.610 1.490 0.945 ;
        RECT 1.115 0.415 1.490 0.610 ;
        RECT 1.115 0.270 1.285 0.415 ;
        RECT 1.850 0.085 2.245 0.580 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__and2b_1

#--------EOF---------

MACRO sky130_fd_sc_hd__and2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.150 0.765 0.450 1.615 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.645 2.200 1.955 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.850 0.785 3.215 1.015 ;
        RECT 0.005 0.105 3.215 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 2.375 1.580 2.680 2.365 ;
        RECT 2.505 0.775 2.680 1.580 ;
        RECT 2.445 0.255 2.680 0.775 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.175 2.015 0.345 2.445 ;
        RECT 0.515 2.185 0.845 2.635 ;
        RECT 0.175 1.785 0.855 2.015 ;
        RECT 0.620 1.135 0.855 1.785 ;
        RECT 1.045 1.475 1.330 2.420 ;
        RECT 1.510 2.165 2.195 2.635 ;
        RECT 2.865 1.680 3.135 2.635 ;
        RECT 1.045 1.325 1.905 1.475 ;
        RECT 1.045 1.305 2.335 1.325 ;
        RECT 0.620 0.805 1.175 1.135 ;
        RECT 1.345 0.945 2.335 1.305 ;
        RECT 0.620 0.655 0.835 0.805 ;
        RECT 0.095 0.085 0.425 0.590 ;
        RECT 0.595 0.280 0.835 0.655 ;
        RECT 1.345 0.610 1.515 0.945 ;
        RECT 1.115 0.415 1.515 0.610 ;
        RECT 1.115 0.270 1.285 0.415 ;
        RECT 1.875 0.085 2.275 0.580 ;
        RECT 2.865 0.085 3.135 0.720 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__and2b_2

#--------EOF---------

MACRO sky130_fd_sc_hd__and2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and2b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.900 1.325 3.155 1.745 ;
        RECT 2.900 0.995 3.205 1.325 ;
        RECT 2.900 0.625 3.155 0.995 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.610 0.995 0.975 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 3.675 1.015 ;
        RECT 0.005 0.105 3.185 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.934000 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.535 2.730 1.745 ;
        RECT 2.440 0.825 2.730 1.535 ;
        RECT 1.525 0.615 2.730 0.825 ;
        RECT 1.525 0.495 1.715 0.615 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.090 2.255 0.425 2.635 ;
        RECT 0.990 2.275 1.320 2.635 ;
        RECT 1.905 2.275 2.235 2.635 ;
        RECT 2.745 2.275 3.075 2.635 ;
        RECT 0.165 1.915 3.505 2.085 ;
        RECT 0.165 1.325 0.335 1.915 ;
        RECT 0.515 1.500 1.315 1.745 ;
        RECT 3.335 1.700 3.505 1.915 ;
        RECT 3.335 1.530 3.545 1.700 ;
        RECT 1.110 1.485 1.315 1.500 ;
        RECT 1.110 1.435 1.320 1.485 ;
        RECT 1.145 1.355 1.320 1.435 ;
        RECT 0.165 0.995 0.425 1.325 ;
        RECT 1.145 0.995 2.260 1.355 ;
        RECT 1.145 0.805 1.355 0.995 ;
        RECT 3.375 0.845 3.545 1.530 ;
        RECT 0.090 0.615 1.355 0.805 ;
        RECT 3.330 0.675 3.545 0.845 ;
        RECT 0.090 0.255 0.425 0.615 ;
        RECT 3.330 0.495 3.500 0.675 ;
        RECT 0.955 0.085 1.285 0.445 ;
        RECT 1.885 0.085 2.215 0.445 ;
        RECT 2.745 0.085 3.075 0.445 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__and2b_4

#--------EOF---------

MACRO sky130_fd_sc_hd__and3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.635 0.635 1.020 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.865 2.125 1.345 2.465 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.145 0.790 1.475 1.215 ;
        RECT 1.145 0.305 1.365 0.790 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.375 0.785 2.295 1.015 ;
        RECT 0.005 0.105 2.295 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 1.940 1.765 2.215 2.465 ;
        RECT 2.045 0.735 2.215 1.765 ;
        RECT 1.955 0.255 2.215 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.085 2.080 0.690 2.635 ;
        RECT 1.515 2.090 1.770 2.635 ;
        RECT 0.085 1.980 0.700 2.080 ;
        RECT 0.515 1.955 0.700 1.980 ;
        RECT 0.085 1.360 0.345 1.810 ;
        RECT 0.515 1.710 0.845 1.955 ;
        RECT 1.015 1.635 1.770 1.885 ;
        RECT 1.000 1.600 1.770 1.635 ;
        RECT 0.985 1.590 1.770 1.600 ;
        RECT 0.980 1.575 1.875 1.590 ;
        RECT 0.960 1.560 1.875 1.575 ;
        RECT 0.940 1.550 1.875 1.560 ;
        RECT 0.915 1.540 1.875 1.550 ;
        RECT 0.845 1.510 1.875 1.540 ;
        RECT 0.825 1.480 1.875 1.510 ;
        RECT 0.805 1.450 1.875 1.480 ;
        RECT 0.775 1.425 1.875 1.450 ;
        RECT 0.740 1.390 1.875 1.425 ;
        RECT 0.710 1.385 1.875 1.390 ;
        RECT 0.710 1.380 1.100 1.385 ;
        RECT 0.710 1.370 1.075 1.380 ;
        RECT 0.710 1.365 1.060 1.370 ;
        RECT 0.710 1.360 1.045 1.365 ;
        RECT 0.085 1.355 1.045 1.360 ;
        RECT 0.085 1.345 1.035 1.355 ;
        RECT 0.085 1.340 1.025 1.345 ;
        RECT 0.085 1.330 1.015 1.340 ;
        RECT 0.085 1.320 1.010 1.330 ;
        RECT 0.085 1.315 1.005 1.320 ;
        RECT 0.085 1.300 0.995 1.315 ;
        RECT 0.085 1.285 0.990 1.300 ;
        RECT 0.085 1.260 0.980 1.285 ;
        RECT 0.085 1.190 0.975 1.260 ;
        RECT 0.805 0.465 0.975 1.190 ;
        RECT 1.645 0.990 1.875 1.385 ;
        RECT 0.085 0.295 0.975 0.465 ;
        RECT 1.535 0.085 1.785 0.625 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__and3_1

#--------EOF---------

MACRO sky130_fd_sc_hd__and3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.470 1.245 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.895 2.125 1.370 2.465 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.750 1.475 1.245 ;
        RECT 1.065 0.305 1.295 0.750 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.345 0.815 2.755 1.015 ;
        RECT 0.020 0.135 2.755 0.815 ;
        RECT 0.145 -0.085 0.315 0.135 ;
        RECT 1.360 0.105 2.755 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 1.970 1.795 2.245 2.465 ;
        RECT 2.075 1.445 2.245 1.795 ;
        RECT 2.060 0.925 2.675 1.445 ;
        RECT 2.060 0.715 2.230 0.925 ;
        RECT 1.980 0.255 2.230 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.085 2.130 0.715 2.635 ;
        RECT 0.100 1.595 0.355 1.960 ;
        RECT 0.525 1.955 0.715 2.130 ;
        RECT 0.525 1.765 0.855 1.955 ;
        RECT 1.080 1.595 1.330 1.890 ;
        RECT 1.555 1.790 1.770 2.635 ;
        RECT 2.415 1.625 2.675 2.635 ;
        RECT 0.100 1.425 1.890 1.595 ;
        RECT 0.640 0.570 0.895 1.425 ;
        RECT 1.660 0.995 1.890 1.425 ;
        RECT 0.105 0.305 0.895 0.570 ;
        RECT 1.475 0.085 1.805 0.580 ;
        RECT 2.400 0.085 2.675 0.745 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__and3_2

#--------EOF---------

MACRO sky130_fd_sc_hd__and3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.115 1.340 0.365 2.335 ;
        RECT 0.115 0.995 0.875 1.340 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.745 1.355 1.340 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 1.900 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER li1 ;
        RECT 2.450 1.760 2.640 2.465 ;
        RECT 3.310 1.765 3.500 2.465 ;
        RECT 3.310 1.760 4.055 1.765 ;
        RECT 2.450 1.535 4.055 1.760 ;
        RECT 3.775 0.845 4.055 1.535 ;
        RECT 2.450 0.615 4.055 0.845 ;
        RECT 2.450 0.515 2.640 0.615 ;
        RECT 3.310 0.255 3.500 0.615 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 0.340 0.105 4.110 1.015 ;
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.545 1.750 0.725 2.465 ;
        RECT 0.895 1.935 1.345 2.635 ;
        RECT 1.520 1.750 1.700 2.465 ;
        RECT 1.910 1.935 2.240 2.635 ;
        RECT 2.810 1.935 3.140 2.635 ;
        RECT 3.670 1.935 4.000 2.635 ;
        RECT 0.545 1.580 2.280 1.750 ;
        RECT 2.070 1.355 2.280 1.580 ;
        RECT 2.070 1.020 3.605 1.355 ;
        RECT 2.070 0.805 2.280 1.020 ;
        RECT 0.465 0.565 0.800 0.805 ;
        RECT 1.535 0.615 2.280 0.805 ;
        RECT 1.535 0.565 1.725 0.615 ;
        RECT 0.465 0.375 1.725 0.565 ;
        RECT 0.465 0.255 0.800 0.375 ;
        RECT 1.905 0.085 2.235 0.445 ;
        RECT 2.810 0.085 3.140 0.445 ;
        RECT 3.670 0.085 4.000 0.445 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__and3_4

#--------EOF---------

MACRO sky130_fd_sc_hd__and3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.955 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.790 2.125 2.265 2.465 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.725 2.395 1.245 ;
        RECT 1.985 0.305 2.185 0.725 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.815 0.935 1.015 ;
        RECT 2.265 0.815 3.215 1.015 ;
        RECT 0.005 0.335 3.215 0.815 ;
        RECT 0.150 0.135 3.215 0.335 ;
        RECT 0.150 -0.085 0.320 0.135 ;
        RECT 2.280 0.105 3.215 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 2.860 1.765 3.135 2.465 ;
        RECT 2.965 0.735 3.135 1.765 ;
        RECT 2.875 0.255 3.135 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 2.125 0.345 2.635 ;
        RECT 0.595 1.245 0.765 2.465 ;
        RECT 1.005 2.130 1.620 2.635 ;
        RECT 1.005 1.595 1.255 1.960 ;
        RECT 1.425 1.955 1.620 2.130 ;
        RECT 2.435 2.090 2.650 2.635 ;
        RECT 1.425 1.765 1.755 1.955 ;
        RECT 1.975 1.595 2.690 1.890 ;
        RECT 1.005 1.425 2.795 1.595 ;
        RECT 0.595 0.995 1.390 1.245 ;
        RECT 0.595 0.905 0.845 0.995 ;
        RECT 0.085 0.085 0.345 0.905 ;
        RECT 0.515 0.485 0.845 0.905 ;
        RECT 1.560 0.570 1.815 1.425 ;
        RECT 2.565 0.995 2.795 1.425 ;
        RECT 1.025 0.305 1.815 0.570 ;
        RECT 2.375 0.085 2.705 0.545 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__and3b_1

#--------EOF---------

MACRO sky130_fd_sc_hd__and3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.745 0.410 1.325 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.815 2.125 2.290 2.465 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.010 0.765 2.420 1.245 ;
        RECT 2.010 0.305 2.220 0.765 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.290 0.815 3.675 1.015 ;
        RECT 0.005 0.135 3.675 0.815 ;
        RECT 0.145 -0.085 0.315 0.135 ;
        RECT 2.305 0.105 3.675 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 2.875 1.795 3.160 2.465 ;
        RECT 2.990 1.445 3.160 1.795 ;
        RECT 2.990 0.925 3.595 1.445 ;
        RECT 2.990 0.715 3.160 0.925 ;
        RECT 2.915 0.255 3.160 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.575 0.400 2.635 ;
        RECT 1.030 2.130 1.645 2.635 ;
        RECT 0.580 1.245 0.855 1.905 ;
        RECT 1.050 1.595 1.285 1.960 ;
        RECT 1.455 1.955 1.645 2.130 ;
        RECT 1.455 1.765 1.785 1.955 ;
        RECT 2.010 1.595 2.200 1.890 ;
        RECT 2.460 1.790 2.675 2.635 ;
        RECT 3.330 1.625 3.595 2.635 ;
        RECT 1.050 1.425 2.820 1.595 ;
        RECT 0.580 1.015 1.415 1.245 ;
        RECT 0.085 0.085 0.355 0.575 ;
        RECT 0.580 0.305 0.855 1.015 ;
        RECT 1.585 0.570 1.840 1.425 ;
        RECT 2.590 0.995 2.820 1.425 ;
        RECT 1.055 0.305 1.840 0.570 ;
        RECT 2.410 0.085 2.740 0.580 ;
        RECT 3.330 0.085 3.595 0.745 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__and3b_2

#--------EOF---------

MACRO sky130_fd_sc_hd__and3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and3b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 3.715 0.615 3.995 1.705 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.020 0.725 1.235 1.340 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 1.715 1.340 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.175 0.335 4.525 1.015 ;
        RECT 0.175 0.105 3.945 0.335 ;
        RECT 0.175 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.934000 ;
    PORT
      LAYER li1 ;
        RECT 2.225 1.535 3.535 1.705 ;
        RECT 3.270 0.845 3.535 1.535 ;
        RECT 2.285 0.615 3.535 0.845 ;
        RECT 2.285 0.515 2.475 0.615 ;
        RECT 3.145 0.255 3.335 0.615 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.730 2.275 1.180 2.635 ;
        RECT 1.745 2.275 2.075 2.635 ;
        RECT 2.645 2.275 2.980 2.635 ;
        RECT 3.505 2.275 3.835 2.635 ;
        RECT 0.150 1.495 0.510 2.165 ;
        RECT 0.680 1.875 4.445 2.105 ;
        RECT 0.150 0.805 0.370 1.495 ;
        RECT 0.680 1.325 0.850 1.875 ;
        RECT 1.280 1.525 2.055 1.695 ;
        RECT 0.540 0.995 0.850 1.325 ;
        RECT 1.885 1.355 2.055 1.525 ;
        RECT 1.885 1.020 3.100 1.355 ;
        RECT 1.885 0.805 2.115 1.020 ;
        RECT 0.150 0.545 0.635 0.805 ;
        RECT 1.420 0.615 2.115 0.805 ;
        RECT 1.420 0.545 1.600 0.615 ;
        RECT 0.150 0.355 1.600 0.545 ;
        RECT 0.150 0.255 0.635 0.355 ;
        RECT 1.780 0.085 2.110 0.445 ;
        RECT 2.645 0.085 2.975 0.445 ;
        RECT 3.505 0.085 3.835 0.445 ;
        RECT 4.165 0.425 4.445 1.875 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__and3b_4

#--------EOF---------

MACRO sky130_fd_sc_hd__and4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.325 2.075 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.885 0.360 1.235 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.415 0.355 1.715 1.325 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.895 0.355 2.175 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.080 0.785 3.215 1.015 ;
        RECT 0.005 0.105 3.215 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 2.795 2.205 3.135 2.465 ;
        RECT 2.875 0.805 3.135 2.205 ;
        RECT 2.795 0.295 3.135 0.805 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.090 2.255 0.425 2.635 ;
        RECT 0.595 1.665 0.845 2.465 ;
        RECT 1.065 1.915 1.395 2.635 ;
        RECT 1.580 1.665 1.830 2.465 ;
        RECT 2.295 1.835 2.625 2.635 ;
        RECT 0.495 1.495 2.685 1.665 ;
        RECT 0.495 0.585 0.665 1.495 ;
        RECT 2.370 1.325 2.685 1.495 ;
        RECT 2.370 1.075 2.700 1.325 ;
        RECT 0.170 0.255 0.665 0.585 ;
        RECT 2.355 0.085 2.625 0.885 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__and4_1

#--------EOF---------

MACRO sky130_fd_sc_hd__and4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.755 0.330 2.075 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.890 0.420 1.245 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.420 1.305 1.590 1.325 ;
        RECT 1.420 0.415 1.720 1.305 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.900 0.415 2.160 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.085 0.785 3.675 1.015 ;
        RECT 0.005 0.105 3.675 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.544500 ;
    PORT
      LAYER li1 ;
        RECT 2.735 1.495 3.070 2.465 ;
        RECT 2.895 0.805 3.070 1.495 ;
        RECT 2.735 0.340 3.070 0.805 ;
        RECT 2.735 0.295 3.065 0.340 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.095 2.255 0.425 2.635 ;
        RECT 0.600 1.665 0.850 2.465 ;
        RECT 1.070 1.915 1.400 2.635 ;
        RECT 1.585 1.665 1.835 2.465 ;
        RECT 2.235 1.835 2.565 2.635 ;
        RECT 3.245 1.835 3.575 2.635 ;
        RECT 0.500 1.495 2.555 1.665 ;
        RECT 0.500 0.585 0.670 1.495 ;
        RECT 2.330 1.315 2.555 1.495 ;
        RECT 2.330 1.075 2.725 1.315 ;
        RECT 0.175 0.255 0.670 0.585 ;
        RECT 2.330 0.085 2.565 0.890 ;
        RECT 3.255 0.085 3.585 0.810 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__and4_2

#--------EOF---------

MACRO sky130_fd_sc_hd__and4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.125 0.765 0.330 1.655 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.840 0.995 1.245 1.325 ;
        RECT 0.890 0.420 1.245 0.995 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.415 0.425 1.700 1.325 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.905 0.935 2.075 1.325 ;
        RECT 1.905 0.730 2.155 0.935 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.135 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 2.535 1.795 2.785 2.465 ;
        RECT 2.615 1.655 2.785 1.795 ;
        RECT 3.375 1.745 3.545 2.465 ;
        RECT 3.375 1.655 4.050 1.745 ;
        RECT 2.615 1.485 4.050 1.655 ;
        RECT 3.800 0.810 4.050 1.485 ;
        RECT 2.535 0.640 4.050 0.810 ;
        RECT 2.535 0.255 2.705 0.640 ;
        RECT 3.375 0.255 3.545 0.640 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.105 1.835 0.385 2.635 ;
        RECT 0.555 1.665 0.765 2.465 ;
        RECT 0.955 1.935 1.285 2.635 ;
        RECT 1.455 1.665 1.645 2.465 ;
        RECT 2.025 1.855 2.355 2.635 ;
        RECT 2.955 1.835 3.205 2.635 ;
        RECT 3.715 1.915 4.045 2.635 ;
        RECT 0.500 1.495 2.415 1.665 ;
        RECT 0.500 0.585 0.670 1.495 ;
        RECT 2.245 1.305 2.415 1.495 ;
        RECT 2.245 1.105 3.585 1.305 ;
        RECT 2.575 1.075 3.585 1.105 ;
        RECT 0.175 0.255 0.670 0.585 ;
        RECT 2.025 0.085 2.335 0.550 ;
        RECT 2.875 0.085 3.205 0.470 ;
        RECT 3.715 0.085 4.045 0.470 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__and4_4

#--------EOF---------

MACRO sky130_fd_sc_hd__and4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.450 1.675 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.520 0.420 1.800 1.695 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.025 0.420 2.295 1.695 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.485 0.665 2.825 1.695 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.745 0.785 3.675 1.015 ;
        RECT 0.005 0.105 3.675 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 3.335 1.495 3.595 2.465 ;
        RECT 3.425 0.805 3.595 1.495 ;
        RECT 3.255 0.340 3.595 0.805 ;
        RECT 3.255 0.295 3.590 0.340 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.170 2.015 0.345 2.465 ;
        RECT 0.515 2.195 0.845 2.635 ;
        RECT 1.150 2.045 1.320 2.465 ;
        RECT 1.555 2.225 2.225 2.635 ;
        RECT 2.440 2.045 2.610 2.465 ;
        RECT 2.810 2.225 3.140 2.635 ;
        RECT 0.170 1.845 0.800 2.015 ;
        RECT 0.630 1.325 0.800 1.845 ;
        RECT 1.150 1.875 3.165 2.045 ;
        RECT 0.630 0.995 0.980 1.325 ;
        RECT 0.630 0.825 0.800 0.995 ;
        RECT 0.170 0.655 0.800 0.825 ;
        RECT 0.170 0.255 0.345 0.655 ;
        RECT 1.150 0.585 1.320 1.875 ;
        RECT 2.995 1.325 3.165 1.875 ;
        RECT 2.995 0.995 3.255 1.325 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.090 0.255 1.320 0.585 ;
        RECT 2.755 0.085 3.085 0.465 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__and4b_1

#--------EOF---------

MACRO sky130_fd_sc_hd__and4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.135 0.740 0.335 1.630 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.420 1.745 1.745 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.960 0.420 2.275 1.695 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.645 2.775 1.615 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.745 0.785 4.135 1.015 ;
        RECT 0.005 0.105 4.135 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.503250 ;
    PORT
      LAYER li1 ;
        RECT 3.340 1.745 3.545 2.465 ;
        RECT 3.340 1.535 4.055 1.745 ;
        RECT 3.425 0.825 4.055 1.535 ;
        RECT 3.260 0.640 4.055 0.825 ;
        RECT 3.260 0.255 3.545 0.640 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.175 2.000 0.345 2.465 ;
        RECT 0.515 2.195 0.845 2.635 ;
        RECT 1.015 2.085 1.185 2.465 ;
        RECT 1.555 2.255 2.225 2.635 ;
        RECT 2.440 2.085 2.610 2.465 ;
        RECT 2.840 2.195 3.170 2.635 ;
        RECT 0.175 1.830 0.805 2.000 ;
        RECT 0.635 1.325 0.805 1.830 ;
        RECT 1.015 1.965 2.610 2.085 ;
        RECT 1.015 1.915 3.165 1.965 ;
        RECT 3.715 1.915 4.050 2.635 ;
        RECT 1.015 1.660 1.315 1.915 ;
        RECT 2.440 1.795 3.165 1.915 ;
        RECT 0.635 0.995 0.975 1.325 ;
        RECT 0.635 0.585 0.805 0.995 ;
        RECT 1.145 0.585 1.315 1.660 ;
        RECT 2.995 1.325 3.165 1.795 ;
        RECT 2.995 0.995 3.255 1.325 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 0.595 0.255 0.805 0.585 ;
        RECT 1.095 0.255 1.315 0.585 ;
        RECT 2.760 0.085 3.090 0.465 ;
        RECT 3.715 0.085 4.050 0.465 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__and4b_2

#--------EOF---------

MACRO sky130_fd_sc_hd__and4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.440 0.765 0.790 1.635 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.815 0.735 4.145 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.345 0.755 3.555 1.325 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.865 0.995 3.085 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.490 0.785 5.055 1.015 ;
        RECT 0.005 0.105 5.055 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.980 1.545 2.160 1.715 ;
        RECT 0.980 0.820 1.260 1.545 ;
        RECT 0.980 0.650 2.080 0.820 ;
        RECT 1.070 0.255 1.240 0.650 ;
        RECT 1.910 0.255 2.080 0.650 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.085 2.085 0.345 2.465 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.410 2.255 1.740 2.635 ;
        RECT 2.250 2.255 2.580 2.635 ;
        RECT 3.475 2.255 3.805 2.635 ;
        RECT 4.635 2.255 4.965 2.635 ;
        RECT 0.085 1.915 4.900 2.085 ;
        RECT 0.085 0.585 0.260 1.915 ;
        RECT 2.380 1.545 4.545 1.715 ;
        RECT 2.380 1.245 2.550 1.545 ;
        RECT 1.440 1.075 2.550 1.245 ;
        RECT 2.380 0.785 2.550 1.075 ;
        RECT 4.730 0.995 4.900 1.915 ;
        RECT 2.380 0.615 2.965 0.785 ;
        RECT 0.085 0.255 0.345 0.585 ;
        RECT 2.795 0.470 2.965 0.615 ;
        RECT 4.390 0.470 4.965 0.810 ;
        RECT 0.570 0.085 0.900 0.470 ;
        RECT 1.410 0.085 1.740 0.470 ;
        RECT 2.285 0.085 2.615 0.445 ;
        RECT 2.795 0.300 4.965 0.470 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
END sky130_fd_sc_hd__and4b_4

#--------EOF---------

MACRO sky130_fd_sc_hd__and4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4bb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.625 0.775 1.955 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.945 1.225 1.115 ;
        RECT 0.605 0.765 0.815 0.945 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.895 1.325 3.080 1.635 ;
        RECT 2.895 0.995 3.125 1.325 ;
        RECT 2.895 0.415 3.080 0.995 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 3.350 1.325 3.545 1.635 ;
        RECT 3.350 0.995 3.605 1.325 ;
        RECT 3.350 0.420 3.545 0.995 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.585 0.785 4.585 1.015 ;
        RECT 0.005 0.695 4.585 0.785 ;
        RECT 0.005 0.335 4.595 0.695 ;
        RECT 0.005 0.105 1.575 0.335 ;
        RECT 3.665 0.145 4.595 0.335 ;
        RECT 3.665 0.105 4.585 0.145 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.425400 ;
    PORT
      LAYER li1 ;
        RECT 4.255 0.255 4.515 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.085 2.135 0.345 2.465 ;
        RECT 0.655 2.255 0.985 2.635 ;
        RECT 0.085 1.455 0.255 2.135 ;
        RECT 1.225 2.085 1.415 2.465 ;
        RECT 1.665 2.255 1.995 2.635 ;
        RECT 2.205 2.085 2.375 2.465 ;
        RECT 2.570 2.255 2.900 2.635 ;
        RECT 3.160 2.085 3.330 2.465 ;
        RECT 3.755 2.255 4.085 2.635 ;
        RECT 1.225 1.915 1.965 2.085 ;
        RECT 1.045 1.575 1.625 1.745 ;
        RECT 1.045 1.455 1.215 1.575 ;
        RECT 0.085 1.285 1.215 1.455 ;
        RECT 1.795 1.405 1.965 1.915 ;
        RECT 0.085 0.585 0.255 1.285 ;
        RECT 1.395 1.235 1.965 1.405 ;
        RECT 2.135 1.915 4.085 2.085 ;
        RECT 1.395 0.755 1.565 1.235 ;
        RECT 2.135 0.925 2.305 1.915 ;
        RECT 0.085 0.255 0.345 0.585 ;
        RECT 0.655 0.085 0.985 0.465 ;
        RECT 1.165 0.425 1.565 0.755 ;
        RECT 1.755 0.595 2.305 0.925 ;
        RECT 2.475 0.425 2.645 1.325 ;
        RECT 3.915 0.995 4.085 1.915 ;
        RECT 1.165 0.255 2.645 0.425 ;
        RECT 3.755 0.085 4.085 0.465 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__and4bb_1

#--------EOF---------

MACRO sky130_fd_sc_hd__and4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4bb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.150 0.995 0.330 1.635 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 3.825 0.765 4.175 1.305 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.910 0.420 3.175 1.275 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 3.350 0.425 3.655 1.405 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.490 0.785 1.830 1.015 ;
        RECT 0.005 0.105 4.595 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.990 1.545 1.320 1.715 ;
        RECT 1.015 0.255 1.240 1.545 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.175 2.055 0.345 2.465 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.490 2.255 2.160 2.635 ;
        RECT 2.395 2.085 2.565 2.465 ;
        RECT 2.735 2.255 3.075 2.635 ;
        RECT 3.245 2.085 3.415 2.465 ;
        RECT 3.755 2.255 4.085 2.635 ;
        RECT 4.255 2.085 4.515 2.465 ;
        RECT 0.175 1.885 1.925 2.055 ;
        RECT 0.500 0.805 0.670 1.885 ;
        RECT 1.755 1.325 1.925 1.885 ;
        RECT 2.235 1.915 3.415 2.085 ;
        RECT 3.585 1.915 4.515 2.085 ;
        RECT 0.175 0.635 0.670 0.805 ;
        RECT 1.415 0.805 1.585 1.325 ;
        RECT 1.755 0.995 2.065 1.325 ;
        RECT 2.235 0.805 2.405 1.915 ;
        RECT 3.585 1.745 3.755 1.915 ;
        RECT 2.575 1.575 3.755 1.745 ;
        RECT 2.575 1.400 2.745 1.575 ;
        RECT 1.415 0.635 2.405 0.805 ;
        RECT 0.175 0.255 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.410 0.085 1.740 0.465 ;
        RECT 2.010 0.255 2.180 0.635 ;
        RECT 4.345 0.585 4.515 1.915 ;
        RECT 3.835 0.085 4.085 0.585 ;
        RECT 4.255 0.255 4.515 0.585 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__and4bb_2

#--------EOF---------

MACRO sky130_fd_sc_hd__and4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__and4bb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 5.485 0.995 5.845 1.620 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.430 0.765 0.780 1.635 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.250 0.755 3.545 1.325 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.680 0.995 3.080 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.490 0.785 4.700 1.015 ;
        RECT 0.005 0.105 5.975 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.960 1.545 2.160 1.715 ;
        RECT 0.960 0.820 1.240 1.545 ;
        RECT 0.960 0.650 2.080 0.820 ;
        RECT 1.070 0.255 1.240 0.650 ;
        RECT 1.910 0.255 2.080 0.650 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.085 2.085 0.345 2.465 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.410 2.255 1.740 2.635 ;
        RECT 2.250 2.255 2.580 2.635 ;
        RECT 3.330 2.255 3.660 2.635 ;
        RECT 4.360 2.255 5.370 2.635 ;
        RECT 5.635 2.085 5.805 2.465 ;
        RECT 0.085 1.915 4.490 2.085 ;
        RECT 0.085 0.585 0.260 1.915 ;
        RECT 2.330 1.545 4.150 1.715 ;
        RECT 2.330 1.245 2.500 1.545 ;
        RECT 4.320 1.325 4.490 1.915 ;
        RECT 1.410 1.075 2.500 1.245 ;
        RECT 2.330 0.785 2.500 1.075 ;
        RECT 3.730 1.155 4.490 1.325 ;
        RECT 4.950 1.915 5.805 2.085 ;
        RECT 3.730 0.995 3.900 1.155 ;
        RECT 4.950 0.825 5.120 1.915 ;
        RECT 2.330 0.615 2.940 0.785 ;
        RECT 0.085 0.255 0.345 0.585 ;
        RECT 2.770 0.470 2.940 0.615 ;
        RECT 4.255 0.470 4.610 0.810 ;
        RECT 4.950 0.655 5.805 0.825 ;
        RECT 0.570 0.085 0.900 0.470 ;
        RECT 1.410 0.085 1.740 0.470 ;
        RECT 2.270 0.085 2.600 0.445 ;
        RECT 2.770 0.300 4.610 0.470 ;
        RECT 4.975 0.085 5.305 0.465 ;
        RECT 5.635 0.255 5.805 0.655 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
END sky130_fd_sc_hd__and4bb_4

#--------EOF---------

MACRO sky130_fd_sc_hd__buf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.985 0.445 1.355 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.375 0.885 ;
        RECT 0.155 -0.085 0.325 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.560 1.295 2.465 ;
        RECT 1.115 0.760 1.295 1.560 ;
        RECT 1.035 0.255 1.295 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.165 1.705 0.345 2.465 ;
        RECT 0.525 1.875 0.855 2.635 ;
        RECT 0.165 1.535 0.840 1.705 ;
        RECT 0.670 1.390 0.840 1.535 ;
        RECT 0.670 1.060 0.945 1.390 ;
        RECT 0.670 0.805 0.840 1.060 ;
        RECT 0.175 0.635 0.840 0.805 ;
        RECT 0.175 0.255 0.345 0.635 ;
        RECT 0.525 0.085 0.855 0.465 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
END sky130_fd_sc_hd__buf_1

#--------EOF---------

MACRO sky130_fd_sc_hd__buf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.440 1.355 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.490 0.785 1.835 1.015 ;
        RECT 0.005 0.105 1.835 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 1.060 1.560 1.315 2.465 ;
        RECT 1.145 0.830 1.315 1.560 ;
        RECT 1.060 0.255 1.315 0.830 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.175 1.705 0.345 2.465 ;
        RECT 0.560 1.875 0.890 2.635 ;
        RECT 0.175 1.535 0.890 1.705 ;
        RECT 0.720 1.325 0.890 1.535 ;
        RECT 1.490 1.485 1.750 2.635 ;
        RECT 0.720 0.995 0.975 1.325 ;
        RECT 0.720 0.805 0.890 0.995 ;
        RECT 0.175 0.635 0.890 0.805 ;
        RECT 0.175 0.255 0.345 0.635 ;
        RECT 0.560 0.085 0.890 0.465 ;
        RECT 1.490 0.085 1.750 0.925 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__buf_2

#--------EOF---------

MACRO sky130_fd_sc_hd__buf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.470 1.315 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.615 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.615 1.185 2.465 ;
        RECT 1.855 1.615 2.025 2.465 ;
        RECT 1.015 1.445 2.025 1.615 ;
        RECT 1.530 0.905 2.025 1.445 ;
        RECT 1.015 0.735 2.025 0.905 ;
        RECT 1.015 0.255 1.185 0.735 ;
        RECT 1.855 0.255 2.025 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.095 1.655 0.425 2.465 ;
        RECT 0.595 1.835 0.835 2.635 ;
        RECT 1.355 1.835 1.685 2.635 ;
        RECT 0.095 1.485 0.810 1.655 ;
        RECT 2.195 1.485 2.525 2.635 ;
        RECT 0.640 1.245 0.810 1.485 ;
        RECT 0.640 1.075 1.140 1.245 ;
        RECT 0.640 0.905 0.810 1.075 ;
        RECT 0.175 0.735 0.810 0.905 ;
        RECT 0.175 0.255 0.345 0.735 ;
        RECT 0.525 0.085 0.765 0.565 ;
        RECT 1.355 0.085 1.685 0.565 ;
        RECT 2.195 0.085 2.525 0.885 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__buf_4

#--------EOF---------

MACRO sky130_fd_sc_hd__buf_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.280 1.075 1.185 1.315 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.265 0.105 4.135 1.015 ;
        RECT 0.265 0.085 0.320 0.105 ;
        RECT 0.150 -0.085 0.320 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER li1 ;
        RECT 1.695 1.615 1.865 2.465 ;
        RECT 2.535 1.615 2.705 2.465 ;
        RECT 3.375 1.615 3.545 2.465 ;
        RECT 1.695 1.445 3.545 1.615 ;
        RECT 2.210 0.905 3.545 1.445 ;
        RECT 1.695 0.735 3.545 0.905 ;
        RECT 1.695 0.255 1.865 0.735 ;
        RECT 2.535 0.255 2.705 0.735 ;
        RECT 3.375 0.255 3.545 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.435 1.485 0.605 2.635 ;
        RECT 0.775 1.655 1.105 2.465 ;
        RECT 1.275 1.835 1.515 2.635 ;
        RECT 2.035 1.835 2.365 2.635 ;
        RECT 2.875 1.835 3.205 2.635 ;
        RECT 0.775 1.485 1.525 1.655 ;
        RECT 3.715 1.485 4.045 2.635 ;
        RECT 1.355 1.245 1.525 1.485 ;
        RECT 1.355 1.075 1.825 1.245 ;
        RECT 1.355 0.905 1.525 1.075 ;
        RECT 0.775 0.735 1.525 0.905 ;
        RECT 0.435 0.085 0.605 0.565 ;
        RECT 0.775 0.255 1.105 0.735 ;
        RECT 1.275 0.085 1.445 0.565 ;
        RECT 2.035 0.085 2.365 0.565 ;
        RECT 2.875 0.085 3.205 0.565 ;
        RECT 3.715 0.085 4.045 0.885 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__buf_6

#--------EOF---------

MACRO sky130_fd_sc_hd__buf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 1.075 1.240 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.135 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 1.855 1.615 2.025 2.465 ;
        RECT 2.695 1.615 2.865 2.465 ;
        RECT 3.535 1.615 3.705 2.465 ;
        RECT 4.375 1.615 4.545 2.465 ;
        RECT 1.855 1.445 4.545 1.615 ;
        RECT 4.290 0.905 4.545 1.445 ;
        RECT 1.855 0.735 4.545 0.905 ;
        RECT 1.855 0.255 2.025 0.735 ;
        RECT 2.695 0.255 2.865 0.735 ;
        RECT 3.535 0.255 3.705 0.735 ;
        RECT 4.375 0.255 4.545 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.095 1.615 0.425 2.465 ;
        RECT 0.595 1.835 0.765 2.635 ;
        RECT 0.935 1.615 1.265 2.465 ;
        RECT 1.435 1.835 1.605 2.635 ;
        RECT 2.195 1.835 2.525 2.635 ;
        RECT 3.035 1.835 3.365 2.635 ;
        RECT 3.875 1.835 4.205 2.635 ;
        RECT 0.095 1.445 1.595 1.615 ;
        RECT 4.715 1.485 5.045 2.635 ;
        RECT 1.420 1.245 1.595 1.445 ;
        RECT 1.420 1.075 4.045 1.245 ;
        RECT 1.420 0.905 1.595 1.075 ;
        RECT 0.175 0.735 1.595 0.905 ;
        RECT 0.175 0.255 0.345 0.735 ;
        RECT 0.515 0.085 0.845 0.565 ;
        RECT 1.015 0.260 1.185 0.735 ;
        RECT 1.355 0.085 1.685 0.565 ;
        RECT 2.195 0.085 2.525 0.565 ;
        RECT 3.035 0.085 3.365 0.565 ;
        RECT 3.875 0.085 4.205 0.565 ;
        RECT 4.715 0.085 5.045 0.885 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__buf_8

#--------EOF---------

MACRO sky130_fd_sc_hd__buf_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.135 1.075 1.660 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.355 1.015 ;
        RECT 0.570 -0.085 0.740 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.615 2.445 2.465 ;
        RECT 3.115 1.615 3.285 2.465 ;
        RECT 3.955 1.615 4.125 2.465 ;
        RECT 4.795 1.615 4.965 2.465 ;
        RECT 5.635 1.615 5.805 2.465 ;
        RECT 6.475 1.615 6.645 2.465 ;
        RECT 2.275 1.445 6.645 1.615 ;
        RECT 4.710 0.905 6.645 1.445 ;
        RECT 2.275 0.735 6.645 0.905 ;
        RECT 2.275 0.255 2.445 0.735 ;
        RECT 3.115 0.255 3.285 0.735 ;
        RECT 3.955 0.255 4.125 0.735 ;
        RECT 4.795 0.255 4.965 0.735 ;
        RECT 5.635 0.255 5.805 0.735 ;
        RECT 6.475 0.255 6.645 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.175 1.835 0.345 2.635 ;
        RECT 0.515 1.615 0.845 2.465 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.355 1.615 1.685 2.465 ;
        RECT 1.855 1.835 2.025 2.635 ;
        RECT 2.615 1.835 2.945 2.635 ;
        RECT 3.455 1.835 3.785 2.635 ;
        RECT 4.295 1.835 4.625 2.635 ;
        RECT 5.135 1.835 5.465 2.635 ;
        RECT 5.975 1.835 6.305 2.635 ;
        RECT 0.515 1.445 2.015 1.615 ;
        RECT 6.815 1.485 7.145 2.635 ;
        RECT 1.840 1.245 2.015 1.445 ;
        RECT 1.840 1.075 4.465 1.245 ;
        RECT 1.840 0.905 2.015 1.075 ;
        RECT 0.595 0.735 2.015 0.905 ;
        RECT 0.095 0.085 0.425 0.565 ;
        RECT 0.595 0.255 0.765 0.735 ;
        RECT 0.935 0.085 1.265 0.565 ;
        RECT 1.435 0.260 1.605 0.735 ;
        RECT 1.775 0.085 2.105 0.565 ;
        RECT 2.615 0.085 2.945 0.565 ;
        RECT 3.455 0.085 3.785 0.565 ;
        RECT 4.295 0.085 4.625 0.565 ;
        RECT 5.135 0.085 5.465 0.565 ;
        RECT 5.975 0.085 6.305 0.565 ;
        RECT 6.815 0.085 7.145 0.885 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
END sky130_fd_sc_hd__buf_12

#--------EOF---------

MACRO sky130_fd_sc_hd__buf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__buf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 2.485 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.755 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER li1 ;
        RECT 3.035 1.615 3.365 2.465 ;
        RECT 3.875 1.615 4.205 2.465 ;
        RECT 4.715 1.615 5.045 2.465 ;
        RECT 5.555 1.615 5.885 2.465 ;
        RECT 6.395 1.615 6.725 2.465 ;
        RECT 7.235 1.615 7.565 2.465 ;
        RECT 8.075 1.615 8.405 2.465 ;
        RECT 8.915 1.615 9.245 2.465 ;
        RECT 9.760 1.615 10.035 2.360 ;
        RECT 3.035 1.445 10.035 1.615 ;
        RECT 9.655 0.905 10.035 1.445 ;
        RECT 3.035 0.735 10.035 0.905 ;
        RECT 3.035 0.260 3.365 0.735 ;
        RECT 3.875 0.260 4.205 0.735 ;
        RECT 4.715 0.260 5.045 0.735 ;
        RECT 5.555 0.260 5.885 0.735 ;
        RECT 6.395 0.260 6.725 0.735 ;
        RECT 7.235 0.260 7.565 0.735 ;
        RECT 8.075 0.260 8.405 0.735 ;
        RECT 8.915 0.260 9.245 0.735 ;
        RECT 9.760 0.365 10.035 0.735 ;
        RECT 3.035 0.255 3.285 0.260 ;
        RECT 3.955 0.255 4.125 0.260 ;
        RECT 4.795 0.255 4.965 0.260 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.175 1.445 0.345 2.635 ;
        RECT 0.515 1.615 0.845 2.465 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.355 1.615 1.685 2.465 ;
        RECT 1.855 1.835 2.025 2.635 ;
        RECT 2.195 1.615 2.525 2.465 ;
        RECT 2.695 1.835 2.865 2.635 ;
        RECT 3.535 1.835 3.705 2.635 ;
        RECT 4.375 1.835 4.545 2.635 ;
        RECT 5.215 1.835 5.385 2.635 ;
        RECT 6.055 1.835 6.225 2.635 ;
        RECT 6.895 1.835 7.065 2.635 ;
        RECT 7.735 1.835 7.905 2.635 ;
        RECT 8.575 1.835 8.745 2.635 ;
        RECT 9.415 1.835 9.585 2.635 ;
        RECT 0.515 1.445 2.865 1.615 ;
        RECT 2.690 1.275 2.865 1.445 ;
        RECT 2.690 1.075 9.410 1.275 ;
        RECT 2.690 0.905 2.865 1.075 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 0.515 0.735 2.865 0.905 ;
        RECT 0.515 0.260 0.845 0.735 ;
        RECT 1.015 0.085 1.185 0.565 ;
        RECT 1.355 0.260 1.685 0.735 ;
        RECT 1.855 0.085 2.025 0.565 ;
        RECT 2.195 0.260 2.525 0.735 ;
        RECT 2.695 0.085 2.865 0.565 ;
        RECT 3.535 0.085 3.705 0.565 ;
        RECT 4.375 0.085 4.545 0.565 ;
        RECT 5.215 0.085 5.385 0.565 ;
        RECT 6.055 0.085 6.225 0.565 ;
        RECT 6.895 0.085 7.065 0.565 ;
        RECT 7.735 0.085 7.905 0.565 ;
        RECT 8.575 0.085 8.745 0.565 ;
        RECT 9.415 0.085 9.585 0.565 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
  END
END sky130_fd_sc_hd__buf_16

#--------EOF---------

MACRO sky130_fd_sc_hd__bufbuf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufbuf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.440 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.490 0.785 6.590 1.015 ;
        RECT 0.005 0.105 6.590 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 3.230 1.615 3.560 2.465 ;
        RECT 4.070 1.615 4.400 2.465 ;
        RECT 4.910 1.615 5.240 2.465 ;
        RECT 5.750 1.615 6.080 2.465 ;
        RECT 3.230 1.445 6.815 1.615 ;
        RECT 6.435 0.905 6.815 1.445 ;
        RECT 3.230 0.735 6.815 0.905 ;
        RECT 3.230 0.260 3.560 0.735 ;
        RECT 4.070 0.260 4.400 0.735 ;
        RECT 4.910 0.260 5.240 0.735 ;
        RECT 5.750 0.260 6.080 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.095 1.615 0.425 2.160 ;
        RECT 0.595 1.785 0.765 2.635 ;
        RECT 0.095 1.445 0.780 1.615 ;
        RECT 1.000 1.545 1.380 2.465 ;
        RECT 0.610 1.325 0.780 1.445 ;
        RECT 0.610 0.995 1.040 1.325 ;
        RECT 1.210 1.275 1.380 1.545 ;
        RECT 1.550 1.615 1.880 2.465 ;
        RECT 2.050 1.785 2.220 2.635 ;
        RECT 2.390 1.615 2.720 2.465 ;
        RECT 2.890 1.785 3.060 2.635 ;
        RECT 3.730 1.835 3.900 2.635 ;
        RECT 4.570 1.835 4.740 2.635 ;
        RECT 5.410 1.835 5.580 2.635 ;
        RECT 6.250 1.835 6.420 2.635 ;
        RECT 1.550 1.445 3.060 1.615 ;
        RECT 2.890 1.275 3.060 1.445 ;
        RECT 1.210 1.075 2.720 1.275 ;
        RECT 2.890 1.075 5.360 1.275 ;
        RECT 0.610 0.905 0.780 0.995 ;
        RECT 0.095 0.735 0.780 0.905 ;
        RECT 1.210 0.825 1.380 1.075 ;
        RECT 2.890 0.905 3.060 1.075 ;
        RECT 0.095 0.260 0.425 0.735 ;
        RECT 0.595 0.085 0.765 0.565 ;
        RECT 1.000 0.260 1.380 0.825 ;
        RECT 1.550 0.735 3.060 0.905 ;
        RECT 1.550 0.260 1.880 0.735 ;
        RECT 2.050 0.085 2.220 0.565 ;
        RECT 2.390 0.260 2.720 0.735 ;
        RECT 2.890 0.085 3.060 0.565 ;
        RECT 3.730 0.085 3.900 0.565 ;
        RECT 4.570 0.085 4.740 0.565 ;
        RECT 5.410 0.085 5.580 0.565 ;
        RECT 6.250 0.085 6.420 0.565 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
  END
END sky130_fd_sc_hd__bufbuf_8

#--------EOF---------

MACRO sky130_fd_sc_hd__bufbuf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufbuf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.960 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.440 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.960 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 11.955 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.150 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.960 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER li1 ;
        RECT 5.235 1.615 5.565 2.465 ;
        RECT 6.075 1.615 6.405 2.465 ;
        RECT 6.915 1.615 7.245 2.465 ;
        RECT 7.755 1.615 8.085 2.465 ;
        RECT 8.595 1.615 8.925 2.465 ;
        RECT 9.435 1.615 9.765 2.465 ;
        RECT 10.275 1.615 10.605 2.465 ;
        RECT 11.115 1.615 11.445 2.465 ;
        RECT 5.235 1.445 11.875 1.615 ;
        RECT 11.620 0.905 11.875 1.445 ;
        RECT 5.235 0.735 11.875 0.905 ;
        RECT 5.235 0.260 5.565 0.735 ;
        RECT 6.075 0.260 6.405 0.735 ;
        RECT 6.915 0.260 7.245 0.735 ;
        RECT 7.755 0.260 8.085 0.735 ;
        RECT 8.595 0.260 8.925 0.735 ;
        RECT 9.435 0.260 9.765 0.735 ;
        RECT 10.275 0.260 10.605 0.735 ;
        RECT 11.115 0.260 11.445 0.735 ;
        RECT 5.235 0.255 5.485 0.260 ;
        RECT 6.155 0.255 6.325 0.260 ;
        RECT 6.995 0.255 7.165 0.260 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.960 2.805 ;
        RECT 0.175 1.445 0.345 2.635 ;
        RECT 0.515 1.445 0.845 2.465 ;
        RECT 1.035 1.615 1.365 2.465 ;
        RECT 1.535 1.785 1.705 2.635 ;
        RECT 1.875 1.615 2.205 2.465 ;
        RECT 2.375 1.785 2.545 2.635 ;
        RECT 2.715 1.615 3.045 2.465 ;
        RECT 3.215 1.835 3.385 2.635 ;
        RECT 3.555 1.615 3.885 2.465 ;
        RECT 4.055 1.835 4.225 2.635 ;
        RECT 4.395 1.615 4.725 2.465 ;
        RECT 4.895 1.835 5.065 2.635 ;
        RECT 5.735 1.835 5.905 2.635 ;
        RECT 6.575 1.835 6.745 2.635 ;
        RECT 7.415 1.835 7.585 2.635 ;
        RECT 8.255 1.835 8.425 2.635 ;
        RECT 9.095 1.835 9.265 2.635 ;
        RECT 9.935 1.835 10.105 2.635 ;
        RECT 10.775 1.835 10.945 2.635 ;
        RECT 11.615 1.835 11.785 2.635 ;
        RECT 1.035 1.445 2.545 1.615 ;
        RECT 2.715 1.445 5.065 1.615 ;
        RECT 0.610 1.275 0.845 1.445 ;
        RECT 2.375 1.275 2.545 1.445 ;
        RECT 4.890 1.275 5.065 1.445 ;
        RECT 0.610 1.075 2.205 1.275 ;
        RECT 2.375 1.075 4.685 1.275 ;
        RECT 4.890 1.075 11.450 1.275 ;
        RECT 0.610 0.905 0.845 1.075 ;
        RECT 2.375 0.905 2.545 1.075 ;
        RECT 4.890 0.905 5.065 1.075 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 0.515 0.260 0.845 0.905 ;
        RECT 1.035 0.735 2.545 0.905 ;
        RECT 2.715 0.735 5.065 0.905 ;
        RECT 1.035 0.260 1.365 0.735 ;
        RECT 1.535 0.085 1.705 0.565 ;
        RECT 1.875 0.260 2.205 0.735 ;
        RECT 2.375 0.085 2.545 0.565 ;
        RECT 2.715 0.260 3.045 0.735 ;
        RECT 3.215 0.085 3.385 0.565 ;
        RECT 3.555 0.260 3.885 0.735 ;
        RECT 4.055 0.085 4.225 0.565 ;
        RECT 4.395 0.260 4.725 0.735 ;
        RECT 4.895 0.085 5.065 0.565 ;
        RECT 5.735 0.085 5.905 0.565 ;
        RECT 6.575 0.085 6.745 0.565 ;
        RECT 7.415 0.085 7.585 0.565 ;
        RECT 8.255 0.085 8.425 0.565 ;
        RECT 9.095 0.085 9.265 0.565 ;
        RECT 9.935 0.085 10.105 0.565 ;
        RECT 10.775 0.085 10.945 0.565 ;
        RECT 11.615 0.085 11.785 0.565 ;
        RECT 0.000 -0.085 11.960 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
  END
END sky130_fd_sc_hd__bufbuf_16

#--------EOF---------

MACRO sky130_fd_sc_hd__bufinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufinv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.505 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.075 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 2.715 1.615 3.045 2.465 ;
        RECT 3.555 1.615 3.885 2.465 ;
        RECT 4.395 1.615 4.725 2.465 ;
        RECT 5.235 1.615 5.565 2.465 ;
        RECT 2.715 1.445 6.355 1.615 ;
        RECT 5.970 0.905 6.355 1.445 ;
        RECT 2.715 0.735 6.355 0.905 ;
        RECT 2.715 0.260 3.045 0.735 ;
        RECT 3.555 0.260 3.885 0.735 ;
        RECT 4.395 0.260 4.725 0.735 ;
        RECT 5.235 0.260 5.565 0.735 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.175 1.445 0.345 2.635 ;
        RECT 0.515 1.545 0.845 2.465 ;
        RECT 0.675 1.275 0.845 1.545 ;
        RECT 1.035 1.615 1.365 2.465 ;
        RECT 1.535 1.785 1.705 2.635 ;
        RECT 1.875 1.615 2.205 2.465 ;
        RECT 2.375 1.785 2.545 2.635 ;
        RECT 3.215 1.835 3.385 2.635 ;
        RECT 4.055 1.835 4.225 2.635 ;
        RECT 4.895 1.835 5.065 2.635 ;
        RECT 5.735 1.835 5.905 2.635 ;
        RECT 1.035 1.445 2.545 1.615 ;
        RECT 2.375 1.275 2.545 1.445 ;
        RECT 0.675 1.075 2.205 1.275 ;
        RECT 2.375 1.075 5.760 1.275 ;
        RECT 0.675 0.905 0.845 1.075 ;
        RECT 2.375 0.905 2.545 1.075 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 0.515 0.260 0.845 0.905 ;
        RECT 1.035 0.735 2.545 0.905 ;
        RECT 1.035 0.260 1.365 0.735 ;
        RECT 1.535 0.085 1.705 0.565 ;
        RECT 1.875 0.260 2.205 0.735 ;
        RECT 2.375 0.085 2.545 0.565 ;
        RECT 3.215 0.085 3.385 0.565 ;
        RECT 4.055 0.085 4.225 0.565 ;
        RECT 4.895 0.085 5.065 0.565 ;
        RECT 5.735 0.085 5.905 0.565 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
END sky130_fd_sc_hd__bufinv_8

#--------EOF---------

MACRO sky130_fd_sc_hd__bufinv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__bufinv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 1.265 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 11.015 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER li1 ;
        RECT 4.295 1.615 4.625 2.465 ;
        RECT 5.135 1.615 5.465 2.465 ;
        RECT 5.975 1.615 6.305 2.465 ;
        RECT 6.815 1.615 7.145 2.465 ;
        RECT 7.655 1.615 7.985 2.465 ;
        RECT 8.495 1.615 8.825 2.465 ;
        RECT 9.335 1.615 9.665 2.465 ;
        RECT 10.175 1.615 10.505 2.465 ;
        RECT 4.295 1.445 10.955 1.615 ;
        RECT 10.680 0.905 10.955 1.445 ;
        RECT 4.295 0.735 10.955 0.905 ;
        RECT 4.295 0.260 4.625 0.735 ;
        RECT 5.135 0.260 5.465 0.735 ;
        RECT 5.975 0.260 6.305 0.735 ;
        RECT 6.815 0.260 7.145 0.735 ;
        RECT 7.655 0.260 7.985 0.735 ;
        RECT 8.495 0.260 8.825 0.735 ;
        RECT 9.335 0.260 9.665 0.735 ;
        RECT 10.175 0.260 10.505 0.735 ;
        RECT 4.295 0.255 4.545 0.260 ;
        RECT 5.215 0.255 5.385 0.260 ;
        RECT 6.055 0.255 6.225 0.260 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.095 1.615 0.425 2.465 ;
        RECT 0.595 1.785 0.765 2.635 ;
        RECT 0.935 1.615 1.265 2.465 ;
        RECT 1.435 1.785 1.605 2.635 ;
        RECT 1.775 1.615 2.105 2.465 ;
        RECT 2.275 1.835 2.445 2.635 ;
        RECT 2.615 1.615 2.945 2.465 ;
        RECT 3.115 1.835 3.285 2.635 ;
        RECT 3.455 1.615 3.785 2.465 ;
        RECT 3.955 1.835 4.125 2.635 ;
        RECT 4.795 1.835 4.965 2.635 ;
        RECT 5.635 1.835 5.805 2.635 ;
        RECT 6.475 1.835 6.645 2.635 ;
        RECT 7.315 1.835 7.485 2.635 ;
        RECT 8.155 1.835 8.325 2.635 ;
        RECT 8.995 1.835 9.165 2.635 ;
        RECT 9.835 1.835 10.005 2.635 ;
        RECT 10.675 1.835 10.845 2.635 ;
        RECT 0.095 1.445 1.605 1.615 ;
        RECT 1.775 1.445 4.125 1.615 ;
        RECT 1.435 1.275 1.605 1.445 ;
        RECT 3.950 1.275 4.125 1.445 ;
        RECT 1.435 1.075 3.745 1.275 ;
        RECT 3.950 1.075 10.510 1.275 ;
        RECT 1.435 0.905 1.605 1.075 ;
        RECT 3.950 0.905 4.125 1.075 ;
        RECT 0.095 0.735 1.605 0.905 ;
        RECT 1.775 0.735 4.125 0.905 ;
        RECT 0.095 0.260 0.425 0.735 ;
        RECT 0.595 0.085 0.765 0.565 ;
        RECT 0.935 0.260 1.265 0.735 ;
        RECT 1.435 0.085 1.605 0.565 ;
        RECT 1.775 0.260 2.105 0.735 ;
        RECT 2.275 0.085 2.445 0.565 ;
        RECT 2.615 0.260 2.945 0.735 ;
        RECT 3.115 0.085 3.285 0.565 ;
        RECT 3.455 0.260 3.785 0.735 ;
        RECT 3.955 0.085 4.125 0.565 ;
        RECT 4.795 0.085 4.965 0.565 ;
        RECT 5.635 0.085 5.805 0.565 ;
        RECT 6.475 0.085 6.645 0.565 ;
        RECT 7.315 0.085 7.485 0.565 ;
        RECT 8.155 0.085 8.325 0.565 ;
        RECT 8.995 0.085 9.165 0.565 ;
        RECT 9.835 0.085 10.005 0.565 ;
        RECT 10.675 0.085 10.845 0.565 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
  END
END sky130_fd_sc_hd__bufinv_16

#--------EOF---------

MACRO sky130_fd_sc_hd__clkbuf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.985 1.275 1.355 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.375 0.885 ;
        RECT 1.065 -0.085 1.235 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.560 0.355 2.465 ;
        RECT 0.085 0.760 0.255 1.560 ;
        RECT 0.085 0.255 0.345 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.525 1.875 0.855 2.635 ;
        RECT 1.035 1.705 1.205 2.465 ;
        RECT 0.540 1.535 1.205 1.705 ;
        RECT 0.540 1.390 0.710 1.535 ;
        RECT 0.425 1.060 0.710 1.390 ;
        RECT 0.540 0.805 0.710 1.060 ;
        RECT 0.540 0.635 1.205 0.805 ;
        RECT 0.525 0.085 0.855 0.465 ;
        RECT 1.035 0.255 1.205 0.635 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
END sky130_fd_sc_hd__clkbuf_1

#--------EOF---------

MACRO sky130_fd_sc_hd__clkbuf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.745 0.785 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.835 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER li1 ;
        RECT 1.060 2.030 1.245 2.435 ;
        RECT 1.060 1.855 1.725 2.030 ;
        RECT 1.385 0.825 1.725 1.855 ;
        RECT 1.040 0.655 1.725 0.825 ;
        RECT 1.040 0.255 1.245 0.655 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.085 1.665 0.355 2.435 ;
        RECT 0.525 1.855 0.855 2.635 ;
        RECT 1.415 2.210 1.750 2.635 ;
        RECT 0.085 1.495 1.215 1.665 ;
        RECT 0.085 0.585 0.255 1.495 ;
        RECT 0.965 0.995 1.215 1.495 ;
        RECT 0.085 0.255 0.345 0.585 ;
        RECT 0.555 0.085 0.830 0.565 ;
        RECT 1.415 0.085 1.750 0.485 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__clkbuf_2

#--------EOF---------

MACRO sky130_fd_sc_hd__clkbuf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.755 0.775 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.745 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER li1 ;
        RECT 1.045 2.005 1.305 2.465 ;
        RECT 1.905 2.005 2.165 2.465 ;
        RECT 1.045 1.835 2.165 2.005 ;
        RECT 1.905 1.585 2.165 1.835 ;
        RECT 1.905 1.415 2.660 1.585 ;
        RECT 2.255 0.905 2.660 1.415 ;
        RECT 1.010 0.735 2.660 0.905 ;
        RECT 1.010 0.345 1.305 0.735 ;
        RECT 1.905 0.345 2.165 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.085 1.665 0.395 2.465 ;
        RECT 0.565 1.835 0.875 2.635 ;
        RECT 1.475 2.175 1.730 2.635 ;
        RECT 2.335 1.765 2.620 2.635 ;
        RECT 0.085 1.495 1.115 1.665 ;
        RECT 0.085 0.585 0.255 1.495 ;
        RECT 0.945 1.245 1.115 1.495 ;
        RECT 0.945 1.075 2.085 1.245 ;
        RECT 0.085 0.255 0.385 0.585 ;
        RECT 0.555 0.085 0.830 0.565 ;
        RECT 1.475 0.085 1.730 0.565 ;
        RECT 2.335 0.085 2.615 0.565 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__clkbuf_4

#--------EOF---------

MACRO sky130_fd_sc_hd__clkbuf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 0.400 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.820 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER li1 ;
        RECT 1.420 1.735 1.680 2.460 ;
        RECT 2.280 1.735 2.540 2.460 ;
        RECT 3.140 1.735 3.400 2.460 ;
        RECT 4.000 1.735 4.260 2.460 ;
        RECT 1.420 1.495 4.730 1.735 ;
        RECT 3.760 0.905 4.730 1.495 ;
        RECT 1.420 0.735 4.730 0.905 ;
        RECT 1.420 0.280 1.680 0.735 ;
        RECT 2.280 0.280 2.540 0.735 ;
        RECT 3.140 0.280 3.400 0.735 ;
        RECT 4.000 0.280 4.260 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.095 1.525 0.390 2.635 ;
        RECT 0.570 1.325 0.820 2.460 ;
        RECT 0.990 1.525 1.250 2.635 ;
        RECT 1.850 1.905 2.110 2.635 ;
        RECT 2.710 1.905 2.970 2.635 ;
        RECT 3.570 1.905 3.830 2.635 ;
        RECT 4.430 1.905 4.725 2.635 ;
        RECT 0.570 1.075 3.590 1.325 ;
        RECT 0.145 0.085 0.390 0.545 ;
        RECT 0.570 0.265 0.820 1.075 ;
        RECT 0.990 0.085 1.250 0.610 ;
        RECT 1.850 0.085 2.110 0.565 ;
        RECT 2.710 0.085 2.970 0.565 ;
        RECT 3.570 0.085 3.830 0.565 ;
        RECT 4.430 0.085 4.730 0.565 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
END sky130_fd_sc_hd__clkbuf_8

#--------EOF---------

MACRO sky130_fd_sc_hd__clkbuf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkbuf_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.400 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.110 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.390 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER li1 ;
        RECT 2.280 1.735 2.540 2.460 ;
        RECT 3.140 1.735 3.400 2.460 ;
        RECT 4.000 1.735 4.260 2.460 ;
        RECT 4.860 1.735 5.120 2.460 ;
        RECT 5.705 1.735 5.965 2.460 ;
        RECT 6.565 1.735 6.825 2.460 ;
        RECT 7.425 1.735 7.685 2.460 ;
        RECT 2.280 1.720 7.685 1.735 ;
        RECT 8.295 1.720 8.585 2.460 ;
        RECT 2.280 1.495 9.025 1.720 ;
        RECT 7.860 0.905 9.025 1.495 ;
        RECT 2.280 0.735 9.025 0.905 ;
        RECT 2.280 0.280 2.540 0.735 ;
        RECT 3.140 0.280 3.400 0.735 ;
        RECT 4.000 0.280 4.260 0.735 ;
        RECT 4.845 0.280 5.120 0.735 ;
        RECT 5.705 0.280 5.965 0.735 ;
        RECT 6.565 0.280 6.825 0.735 ;
        RECT 7.425 0.280 7.685 0.735 ;
        RECT 8.295 0.280 8.555 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.095 1.825 0.390 2.635 ;
        RECT 0.570 1.325 0.815 2.465 ;
        RECT 0.990 1.825 1.250 2.635 ;
        RECT 1.850 2.630 8.125 2.635 ;
        RECT 1.430 1.325 1.680 2.460 ;
        RECT 1.850 1.835 2.110 2.630 ;
        RECT 2.710 1.905 2.970 2.630 ;
        RECT 3.570 1.905 3.830 2.630 ;
        RECT 4.430 1.905 4.690 2.630 ;
        RECT 5.290 1.905 5.535 2.630 ;
        RECT 6.150 1.905 6.395 2.630 ;
        RECT 7.010 1.905 7.255 2.630 ;
        RECT 7.870 1.905 8.125 2.630 ;
        RECT 8.755 1.890 9.025 2.635 ;
        RECT 0.570 1.075 7.690 1.325 ;
        RECT 0.085 0.085 0.390 0.595 ;
        RECT 0.570 0.265 0.820 1.075 ;
        RECT 0.990 0.085 1.250 0.610 ;
        RECT 1.430 0.265 1.680 1.075 ;
        RECT 1.850 0.085 2.110 0.645 ;
        RECT 2.710 0.085 2.970 0.565 ;
        RECT 3.570 0.085 3.830 0.565 ;
        RECT 4.430 0.085 4.675 0.565 ;
        RECT 5.290 0.085 5.535 0.565 ;
        RECT 6.145 0.085 6.395 0.565 ;
        RECT 7.005 0.085 7.255 0.565 ;
        RECT 7.865 0.085 8.125 0.565 ;
        RECT 8.725 0.085 9.025 0.565 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
  END
END sky130_fd_sc_hd__clkbuf_16

#--------EOF---------

MACRO sky130_fd_sc_hd__clkdlybuf4s15_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s15_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.560 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.495 0.785 3.115 1.015 ;
        RECT 0.005 0.105 3.640 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.376300 ;
    PORT
      LAYER li1 ;
        RECT 3.210 1.760 3.595 2.465 ;
        RECT 3.365 0.545 3.595 1.760 ;
        RECT 3.210 0.285 3.595 0.545 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.665 0.425 2.465 ;
        RECT 0.595 1.835 0.925 2.635 ;
        RECT 1.385 1.835 1.760 2.465 ;
        RECT 0.085 1.495 1.215 1.665 ;
        RECT 0.730 0.885 1.215 1.495 ;
        RECT 0.085 0.715 1.215 0.885 ;
        RECT 1.590 1.250 1.760 1.835 ;
        RECT 1.930 1.590 2.410 2.465 ;
        RECT 2.640 1.760 3.040 2.635 ;
        RECT 1.930 1.420 3.195 1.590 ;
        RECT 1.590 1.055 2.685 1.250 ;
        RECT 1.590 0.825 1.760 1.055 ;
        RECT 2.855 0.885 3.195 1.420 ;
        RECT 0.085 0.255 0.425 0.715 ;
        RECT 0.595 0.085 0.910 0.545 ;
        RECT 1.385 0.255 1.760 0.825 ;
        RECT 1.930 0.715 3.195 0.885 ;
        RECT 1.930 0.255 2.260 0.715 ;
        RECT 2.710 0.085 3.040 0.545 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s15_1

#--------EOF---------

MACRO sky130_fd_sc_hd__clkdlybuf4s15_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s15_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.060 0.555 1.625 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.535 0.785 2.620 1.015 ;
        RECT 0.005 0.105 4.135 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.397600 ;
    PORT
      LAYER li1 ;
        RECT 3.070 1.485 3.550 2.465 ;
        RECT 3.355 0.640 3.550 1.485 ;
        RECT 3.050 0.255 3.550 0.640 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 1.965 0.430 2.465 ;
        RECT 0.600 2.135 0.930 2.635 ;
        RECT 0.085 1.795 1.060 1.965 ;
        RECT 0.890 1.245 1.060 1.795 ;
        RECT 1.230 1.785 1.660 2.465 ;
        RECT 1.830 1.965 2.100 2.465 ;
        RECT 2.550 2.135 2.880 2.635 ;
        RECT 1.830 1.790 2.900 1.965 ;
        RECT 1.490 1.485 1.660 1.785 ;
        RECT 0.890 1.075 1.320 1.245 ;
        RECT 1.490 1.075 2.415 1.485 ;
        RECT 2.730 1.245 2.900 1.790 ;
        RECT 3.720 1.485 4.055 2.635 ;
        RECT 2.730 1.075 3.185 1.245 ;
        RECT 0.890 0.890 1.060 1.075 ;
        RECT 1.490 0.905 1.660 1.075 ;
        RECT 2.730 0.905 2.900 1.075 ;
        RECT 0.085 0.720 1.060 0.890 ;
        RECT 0.085 0.255 0.415 0.720 ;
        RECT 0.585 0.085 0.915 0.550 ;
        RECT 1.280 0.255 1.660 0.905 ;
        RECT 1.830 0.735 2.900 0.905 ;
        RECT 1.830 0.255 2.100 0.735 ;
        RECT 2.550 0.085 2.880 0.565 ;
        RECT 3.720 0.085 4.055 0.645 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s15_2

#--------EOF---------

MACRO sky130_fd_sc_hd__clkdlybuf4s18_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s18_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.055 0.550 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.530 0.785 3.115 1.015 ;
        RECT 0.005 0.105 3.640 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.376300 ;
    PORT
      LAYER li1 ;
        RECT 3.220 1.760 3.590 2.465 ;
        RECT 3.365 0.545 3.590 1.760 ;
        RECT 3.210 0.255 3.590 0.545 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.095 1.665 0.425 2.465 ;
        RECT 0.595 1.835 0.925 2.635 ;
        RECT 1.385 1.835 1.760 2.465 ;
        RECT 0.095 1.495 1.215 1.665 ;
        RECT 0.720 0.885 1.215 1.495 ;
        RECT 0.095 0.715 1.215 0.885 ;
        RECT 1.590 1.250 1.760 1.835 ;
        RECT 1.930 1.590 2.260 2.465 ;
        RECT 2.710 1.760 3.040 2.635 ;
        RECT 1.930 1.420 3.195 1.590 ;
        RECT 1.590 1.055 2.685 1.250 ;
        RECT 1.590 0.825 1.760 1.055 ;
        RECT 2.855 0.885 3.195 1.420 ;
        RECT 0.095 0.255 0.425 0.715 ;
        RECT 0.595 0.085 0.910 0.545 ;
        RECT 1.385 0.255 1.760 0.825 ;
        RECT 1.930 0.715 3.195 0.885 ;
        RECT 1.930 0.255 2.260 0.715 ;
        RECT 2.710 0.085 3.040 0.545 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s18_1

#--------EOF---------

MACRO sky130_fd_sc_hd__clkdlybuf4s18_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s18_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.560 1.290 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.535 0.785 2.635 1.015 ;
        RECT 0.005 0.105 3.675 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.397600 ;
    PORT
      LAYER li1 ;
        RECT 2.715 1.525 3.150 2.465 ;
        RECT 2.715 1.420 3.180 1.525 ;
        RECT 3.010 0.945 3.180 1.420 ;
        RECT 2.965 0.780 3.180 0.945 ;
        RECT 2.965 0.640 3.150 0.780 ;
        RECT 2.705 0.270 3.150 0.640 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.630 0.430 2.465 ;
        RECT 0.600 1.800 0.930 2.635 ;
        RECT 1.110 1.800 1.440 2.465 ;
        RECT 0.085 1.460 1.055 1.630 ;
        RECT 0.730 0.905 1.055 1.460 ;
        RECT 0.085 0.735 1.055 0.905 ;
        RECT 1.270 1.255 1.440 1.800 ;
        RECT 1.630 1.630 1.960 2.465 ;
        RECT 2.130 1.800 2.545 2.635 ;
        RECT 1.630 1.460 2.545 1.630 ;
        RECT 3.320 1.625 3.595 2.635 ;
        RECT 1.270 1.075 2.205 1.255 ;
        RECT 2.375 1.245 2.545 1.460 ;
        RECT 2.375 1.075 2.840 1.245 ;
        RECT 0.085 0.270 0.415 0.735 ;
        RECT 1.270 0.600 1.440 1.075 ;
        RECT 2.375 0.905 2.545 1.075 ;
        RECT 0.585 0.085 0.915 0.565 ;
        RECT 1.160 0.270 1.440 0.600 ;
        RECT 1.630 0.735 2.545 0.905 ;
        RECT 1.630 0.270 1.960 0.735 ;
        RECT 2.165 0.085 2.535 0.565 ;
        RECT 3.320 0.085 3.595 0.645 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s18_2

#--------EOF---------

MACRO sky130_fd_sc_hd__clkdlybuf4s25_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s25_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.485 1.320 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.530 0.785 2.920 1.015 ;
        RECT 0.005 0.105 3.675 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.702900 ;
    PORT
      LAYER li1 ;
        RECT 3.035 1.565 3.595 2.465 ;
        RECT 3.230 0.640 3.595 1.565 ;
        RECT 3.015 0.255 3.595 0.640 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.660 0.430 2.465 ;
        RECT 0.600 1.830 0.925 2.635 ;
        RECT 1.195 1.790 1.645 2.465 ;
        RECT 0.085 1.490 1.005 1.660 ;
        RECT 0.655 1.295 1.005 1.490 ;
        RECT 0.655 1.025 1.105 1.295 ;
        RECT 1.470 1.250 1.645 1.790 ;
        RECT 1.815 1.665 2.065 2.465 ;
        RECT 2.235 1.835 2.845 2.635 ;
        RECT 1.815 1.495 2.765 1.665 ;
        RECT 2.595 1.325 2.765 1.495 ;
        RECT 1.470 1.075 2.420 1.250 ;
        RECT 0.655 0.905 1.005 1.025 ;
        RECT 0.085 0.735 1.005 0.905 ;
        RECT 1.470 0.855 1.645 1.075 ;
        RECT 2.595 0.990 3.050 1.325 ;
        RECT 2.595 0.905 2.765 0.990 ;
        RECT 0.085 0.255 0.410 0.735 ;
        RECT 0.580 0.085 0.910 0.565 ;
        RECT 1.175 0.255 1.645 0.855 ;
        RECT 1.815 0.735 2.765 0.905 ;
        RECT 1.815 0.255 2.065 0.735 ;
        RECT 2.240 0.085 2.845 0.565 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s25_1

#--------EOF---------

MACRO sky130_fd_sc_hd__clkdlybuf4s25_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s25_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.495 1.615 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.495 0.785 2.545 1.015 ;
        RECT 0.005 0.105 3.605 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.497000 ;
    PORT
      LAYER li1 ;
        RECT 2.770 1.625 3.095 2.460 ;
        RECT 2.865 1.275 3.095 1.625 ;
        RECT 2.865 0.765 3.595 1.275 ;
        RECT 2.865 0.615 3.095 0.765 ;
        RECT 2.770 0.285 3.095 0.615 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.095 1.955 0.345 2.465 ;
        RECT 0.575 2.125 0.905 2.635 ;
        RECT 0.095 1.785 0.835 1.955 ;
        RECT 0.665 1.750 0.835 1.785 ;
        RECT 0.665 1.325 1.005 1.750 ;
        RECT 1.175 1.425 1.440 2.465 ;
        RECT 1.695 1.745 1.945 2.465 ;
        RECT 2.135 1.915 2.465 2.635 ;
        RECT 1.695 1.500 2.595 1.745 ;
        RECT 3.265 1.635 3.595 2.635 ;
        RECT 1.205 1.325 1.440 1.425 ;
        RECT 0.665 0.995 1.035 1.325 ;
        RECT 1.205 0.995 2.165 1.325 ;
        RECT 0.665 0.810 0.840 0.995 ;
        RECT 0.095 0.640 0.840 0.810 ;
        RECT 1.205 0.780 1.425 0.995 ;
        RECT 2.335 0.805 2.595 1.500 ;
        RECT 0.095 0.305 0.345 0.640 ;
        RECT 0.575 0.085 0.905 0.470 ;
        RECT 1.095 0.255 1.425 0.780 ;
        RECT 1.615 0.635 2.595 0.805 ;
        RECT 1.615 0.255 1.945 0.635 ;
        RECT 2.135 0.085 2.465 0.465 ;
        RECT 3.265 0.085 3.595 0.550 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s25_2

#--------EOF---------

MACRO sky130_fd_sc_hd__clkdlybuf4s50_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s50_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.535 1.290 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.535 0.785 3.095 1.015 ;
        RECT 0.005 0.105 3.675 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504100 ;
    PORT
      LAYER li1 ;
        RECT 3.190 1.690 3.595 2.465 ;
        RECT 3.345 0.640 3.595 1.690 ;
        RECT 3.190 0.255 3.595 0.640 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.630 0.430 2.465 ;
        RECT 0.600 1.800 0.930 2.635 ;
        RECT 0.085 1.460 1.055 1.630 ;
        RECT 0.705 1.315 1.055 1.460 ;
        RECT 1.380 1.320 1.730 2.465 ;
        RECT 1.990 1.665 2.240 2.465 ;
        RECT 2.690 1.835 3.020 2.635 ;
        RECT 1.990 1.495 2.580 1.665 ;
        RECT 2.410 1.325 2.580 1.495 ;
        RECT 0.705 1.025 1.135 1.315 ;
        RECT 1.380 1.070 2.240 1.320 ;
        RECT 0.705 0.905 1.055 1.025 ;
        RECT 0.085 0.735 1.055 0.905 ;
        RECT 0.085 0.255 0.415 0.735 ;
        RECT 0.585 0.085 0.915 0.565 ;
        RECT 1.380 0.255 1.730 1.070 ;
        RECT 2.410 0.995 3.175 1.325 ;
        RECT 2.410 0.900 2.580 0.995 ;
        RECT 1.990 0.730 2.580 0.900 ;
        RECT 1.990 0.255 2.240 0.730 ;
        RECT 2.690 0.085 3.020 0.600 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s50_1

#--------EOF---------

MACRO sky130_fd_sc_hd__clkdlybuf4s50_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkdlybuf4s50_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.480 1.285 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.535 0.785 3.090 1.015 ;
        RECT 0.005 0.105 4.135 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.390500 ;
    PORT
      LAYER li1 ;
        RECT 3.185 1.530 3.625 2.465 ;
        RECT 3.345 0.640 3.625 1.530 ;
        RECT 3.185 0.270 3.625 0.640 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 1.630 0.430 2.465 ;
        RECT 0.600 1.800 0.930 2.635 ;
        RECT 1.390 1.785 1.795 2.465 ;
        RECT 0.085 1.455 1.270 1.630 ;
        RECT 0.850 1.245 1.270 1.455 ;
        RECT 1.625 1.245 1.795 1.785 ;
        RECT 1.985 1.630 2.235 2.465 ;
        RECT 2.685 1.800 3.015 2.635 ;
        RECT 3.795 1.800 4.055 2.635 ;
        RECT 1.985 1.460 2.645 1.630 ;
        RECT 2.475 1.325 2.645 1.460 ;
        RECT 0.765 1.075 1.435 1.245 ;
        RECT 1.625 1.075 2.305 1.245 ;
        RECT 0.850 0.905 1.270 1.075 ;
        RECT 0.085 0.735 1.270 0.905 ;
        RECT 1.625 0.900 1.795 1.075 ;
        RECT 2.475 0.995 3.175 1.325 ;
        RECT 2.475 0.905 2.645 0.995 ;
        RECT 0.085 0.270 0.415 0.735 ;
        RECT 0.585 0.085 0.915 0.565 ;
        RECT 1.440 0.270 1.795 0.900 ;
        RECT 1.985 0.735 2.645 0.905 ;
        RECT 1.985 0.270 2.235 0.735 ;
        RECT 2.685 0.085 3.015 0.565 ;
        RECT 3.795 0.085 4.055 0.635 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__clkdlybuf4s50_2

#--------EOF---------

MACRO sky130_fd_sc_hd__clkinv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.315000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.375 0.325 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.290 0.845 2.465 ;
        RECT 0.515 0.760 1.295 1.290 ;
        RECT 0.515 0.255 0.840 0.760 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 0.420 0.105 1.375 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.085 1.665 0.345 2.635 ;
        RECT 1.015 1.665 1.295 2.635 ;
        RECT 1.010 0.085 1.295 0.590 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
END sky130_fd_sc_hd__clkinv_1

#--------EOF---------

MACRO sky130_fd_sc_hd__clkinv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.576000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.065 1.305 1.290 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.662600 ;
    PORT
      LAYER li1 ;
        RECT 0.155 1.630 0.410 2.435 ;
        RECT 1.010 1.630 1.270 2.435 ;
        RECT 0.155 1.460 1.755 1.630 ;
        RECT 1.475 0.895 1.755 1.460 ;
        RECT 1.025 0.725 1.755 0.895 ;
        RECT 1.025 0.280 1.250 0.725 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 0.470 0.105 1.835 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.580 1.800 0.840 2.635 ;
        RECT 1.440 1.800 1.695 2.635 ;
        RECT 0.560 0.085 0.855 0.610 ;
        RECT 1.420 0.085 1.750 0.555 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__clkinv_2

#--------EOF---------

MACRO sky130_fd_sc_hd__clkinv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.065 2.660 1.290 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.075200 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.630 0.860 2.435 ;
        RECT 1.465 1.630 1.720 2.435 ;
        RECT 2.320 1.630 2.580 2.435 ;
        RECT 0.105 1.460 3.135 1.630 ;
        RECT 0.105 0.895 0.275 1.460 ;
        RECT 2.835 0.895 3.135 1.460 ;
        RECT 0.105 0.725 3.135 0.895 ;
        RECT 1.030 0.280 1.290 0.725 ;
        RECT 1.890 0.280 2.145 0.725 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 0.410 0.105 2.835 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.800 0.430 2.635 ;
        RECT 1.030 1.800 1.290 2.635 ;
        RECT 1.890 1.800 2.150 2.635 ;
        RECT 2.750 1.800 3.135 2.635 ;
        RECT 0.565 0.085 0.860 0.555 ;
        RECT 1.460 0.085 1.720 0.555 ;
        RECT 2.315 0.085 2.615 0.555 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__clkinv_4

#--------EOF---------

MACRO sky130_fd_sc_hd__clkinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.304000 ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.035 4.865 1.290 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150 -0.085 0.320 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.090400 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.630 0.805 2.435 ;
        RECT 1.405 1.630 1.645 2.435 ;
        RECT 2.245 1.630 2.495 2.435 ;
        RECT 3.080 1.630 3.325 2.435 ;
        RECT 3.920 1.630 4.175 2.435 ;
        RECT 4.765 1.630 5.005 2.435 ;
        RECT 0.115 1.460 5.440 1.630 ;
        RECT 0.115 0.865 0.285 1.460 ;
        RECT 5.170 0.865 5.440 1.460 ;
        RECT 0.115 0.695 5.440 0.865 ;
        RECT 1.535 0.280 1.725 0.695 ;
        RECT 2.395 0.280 2.585 0.695 ;
        RECT 3.255 0.280 3.445 0.695 ;
        RECT 4.115 0.280 4.305 0.695 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 0.945 0.105 4.895 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.135 1.800 0.395 2.635 ;
        RECT 0.975 1.800 1.235 2.635 ;
        RECT 1.815 1.800 2.075 2.635 ;
        RECT 2.665 1.800 2.910 2.635 ;
        RECT 3.495 1.800 3.750 2.635 ;
        RECT 4.345 1.800 4.595 2.635 ;
        RECT 5.175 1.800 5.430 2.635 ;
        RECT 1.035 0.085 1.365 0.525 ;
        RECT 1.895 0.085 2.225 0.525 ;
        RECT 2.755 0.085 3.085 0.525 ;
        RECT 3.615 0.085 3.945 0.525 ;
        RECT 4.475 0.085 4.805 0.525 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
END sky130_fd_sc_hd__clkinv_8

#--------EOF---------

MACRO sky130_fd_sc_hd__clkinv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.608000 ;
    PORT
      LAYER met1 ;
        RECT 1.465 1.260 2.215 1.305 ;
        RECT 9.285 1.260 10.035 1.305 ;
        RECT 1.465 1.120 10.035 1.260 ;
        RECT 1.465 1.075 2.215 1.120 ;
        RECT 9.285 1.075 10.035 1.120 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER li1 ;
        RECT 0.575 1.665 0.830 2.465 ;
        RECT 1.435 1.665 1.690 2.450 ;
        RECT 2.325 1.665 2.550 2.465 ;
        RECT 3.155 1.665 3.410 2.450 ;
        RECT 4.015 1.665 4.255 2.450 ;
        RECT 4.905 1.665 5.280 2.450 ;
        RECT 5.925 1.665 6.175 2.450 ;
        RECT 6.785 1.665 7.035 2.450 ;
        RECT 7.645 1.665 7.895 2.450 ;
        RECT 8.505 1.665 8.755 2.450 ;
        RECT 9.365 1.665 9.605 2.450 ;
        RECT 10.225 1.665 10.480 2.450 ;
        RECT 0.575 1.455 10.480 1.665 ;
        RECT 2.325 1.415 8.755 1.455 ;
        RECT 2.325 0.280 2.550 1.415 ;
        RECT 3.155 0.280 3.410 1.415 ;
        RECT 4.015 0.280 4.255 1.415 ;
        RECT 4.905 0.280 5.255 1.415 ;
        RECT 5.925 0.280 6.175 1.415 ;
        RECT 6.785 0.280 7.035 1.415 ;
        RECT 7.645 0.280 7.895 1.415 ;
        RECT 8.505 0.280 8.755 1.415 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 1.735 0.105 9.315 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.140 1.495 0.405 2.635 ;
        RECT 1.000 1.835 1.260 2.635 ;
        RECT 1.865 1.835 2.120 2.635 ;
        RECT 2.720 1.835 2.980 2.635 ;
        RECT 3.585 1.835 3.840 2.635 ;
        RECT 4.465 1.835 4.720 2.635 ;
        RECT 5.490 2.120 5.750 2.635 ;
        RECT 5.490 1.835 5.745 2.120 ;
        RECT 6.355 1.835 6.610 2.635 ;
        RECT 7.215 1.835 7.470 2.635 ;
        RECT 8.075 1.835 8.330 2.635 ;
        RECT 8.935 1.835 9.190 2.635 ;
        RECT 9.795 1.835 10.050 2.635 ;
        RECT 10.650 1.835 10.910 2.635 ;
        RECT 0.345 0.895 2.155 1.275 ;
        RECT 8.930 0.895 10.710 1.275 ;
        RECT 1.855 0.085 2.125 0.610 ;
        RECT 2.720 0.085 2.985 0.610 ;
        RECT 3.580 0.085 3.845 0.610 ;
        RECT 4.465 0.085 4.730 0.610 ;
        RECT 5.490 0.085 5.755 0.610 ;
        RECT 6.350 0.085 6.575 0.610 ;
        RECT 7.210 0.085 7.475 0.610 ;
        RECT 8.070 0.085 8.335 0.610 ;
        RECT 8.930 0.085 9.195 0.610 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 1.525 1.105 1.695 1.275 ;
        RECT 1.985 1.105 2.155 1.275 ;
        RECT 9.345 1.105 9.515 1.275 ;
        RECT 9.805 1.105 9.975 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
  END
END sky130_fd_sc_hd__clkinv_16

#--------EOF---------

MACRO sky130_fd_sc_hd__clkinvlp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinvlp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.665000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.995 0.600 1.665 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.185 0.205 1.555 1.015 ;
        RECT 0.185 0.085 0.315 0.205 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.436750 ;
    PORT
      LAYER li1 ;
        RECT 0.810 0.750 1.235 2.455 ;
        RECT 0.810 0.315 1.445 0.750 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.225 2.625 1.740 2.635 ;
        RECT 0.225 1.835 0.555 2.625 ;
        RECT 1.440 1.455 1.740 2.625 ;
        RECT 0.295 0.085 0.625 0.745 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__clkinvlp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__clkinvlp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__clkinvlp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.330000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.745 0.425 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.095 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.714000 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.295 0.955 2.465 ;
        RECT 1.685 1.295 2.015 2.465 ;
        RECT 0.595 1.015 2.015 1.295 ;
        RECT 0.595 0.680 0.955 1.015 ;
        RECT 0.595 0.255 1.215 0.680 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.095 1.495 0.425 2.635 ;
        RECT 1.155 1.465 1.485 2.635 ;
        RECT 2.215 1.465 2.545 2.635 ;
        RECT 0.095 0.085 0.425 0.575 ;
        RECT 1.675 0.085 2.005 0.775 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__clkinvlp_4

#--------EOF---------

MACRO sky130_fd_sc_hd__conb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__conb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.605 1.740 ;
    END
  END HI
  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.775 0.915 1.295 2.465 ;
    END
  END LO
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.275 1.910 0.605 2.635 ;
        RECT 0.775 0.085 1.115 0.745 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
END sky130_fd_sc_hd__conb_1

#--------EOF---------

MACRO sky130_fd_sc_hd__decap_3
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__decap_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.375 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.085 1.545 1.295 2.635 ;
        RECT 0.085 0.835 0.605 1.375 ;
        RECT 0.775 1.005 1.295 1.545 ;
        RECT 0.085 0.085 1.295 0.835 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
END sky130_fd_sc_hd__decap_3

#--------EOF---------

MACRO sky130_fd_sc_hd__decap_4
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__decap_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.835 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.085 1.545 1.755 2.635 ;
        RECT 0.085 0.855 0.835 1.375 ;
        RECT 1.005 1.025 1.755 1.545 ;
        RECT 0.085 0.085 1.755 0.855 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__decap_4

#--------EOF---------

MACRO sky130_fd_sc_hd__decap_6
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__decap_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.755 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.085 1.545 2.675 2.635 ;
        RECT 0.085 0.855 1.295 1.375 ;
        RECT 1.465 1.025 2.675 1.545 ;
        RECT 0.085 0.085 2.675 0.855 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__decap_6

#--------EOF---------

MACRO sky130_fd_sc_hd__decap_8
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__decap_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.675 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.545 3.595 2.635 ;
        RECT 0.085 0.855 1.735 1.375 ;
        RECT 1.905 1.025 3.595 1.545 ;
        RECT 0.085 0.085 3.595 0.855 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__decap_8

#--------EOF---------

MACRO sky130_fd_sc_hd__decap_12
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__decap_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.515 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.085 1.545 5.430 2.635 ;
        RECT 0.085 0.855 2.665 1.375 ;
        RECT 2.835 1.025 5.430 1.545 ;
        RECT 0.085 0.085 5.430 0.855 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__decap_12

#--------EOF---------

MACRO sky130_fd_sc_hd__dfbbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfbbn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.960 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK_N
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.745 1.005 2.155 1.625 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 9.235 1.095 9.690 1.325 ;
    END
  END RESET_B
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 3.765 0.920 4.055 0.965 ;
        RECT 7.515 0.920 7.805 0.965 ;
        RECT 3.765 0.780 7.805 0.920 ;
        RECT 3.765 0.735 4.055 0.780 ;
        RECT 7.515 0.735 7.805 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.960 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 9.620 1.005 11.955 1.015 ;
        RECT 3.900 0.785 6.175 1.005 ;
        RECT 7.785 0.785 11.955 1.005 ;
        RECT 0.005 0.105 11.955 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.150 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.960 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 11.615 1.455 11.875 2.465 ;
        RECT 11.665 0.825 11.875 1.455 ;
        RECT 11.615 0.255 11.875 0.825 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 10.200 1.630 10.485 2.465 ;
        RECT 10.305 0.715 10.485 1.630 ;
        RECT 10.200 0.255 10.485 0.715 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.960 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.175 0.635 0.840 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.235 2.465 ;
        RECT 1.430 2.135 1.785 2.635 ;
        RECT 1.955 1.965 2.125 2.465 ;
        RECT 2.335 2.250 3.165 2.420 ;
        RECT 1.405 1.795 2.125 1.965 ;
        RECT 1.405 0.825 1.575 1.795 ;
        RECT 2.325 1.575 2.825 1.955 ;
        RECT 1.405 0.635 2.125 0.825 ;
        RECT 2.325 0.705 2.545 1.575 ;
        RECT 2.995 1.405 3.165 2.250 ;
        RECT 3.405 2.205 3.785 2.635 ;
        RECT 4.085 2.035 4.255 2.375 ;
        RECT 3.335 1.785 4.685 2.035 ;
        RECT 4.875 1.915 5.205 2.635 ;
        RECT 6.250 2.250 7.080 2.420 ;
        RECT 7.320 2.255 7.700 2.635 ;
        RECT 3.335 1.575 3.585 1.785 ;
        RECT 4.095 1.405 4.345 1.485 ;
        RECT 2.995 1.235 4.345 1.405 ;
        RECT 2.995 1.195 3.415 1.235 ;
        RECT 2.725 0.645 3.075 1.015 ;
        RECT 1.430 0.085 1.785 0.465 ;
        RECT 1.955 0.305 2.125 0.635 ;
        RECT 3.245 0.465 3.415 1.195 ;
        RECT 4.125 1.155 4.345 1.235 ;
        RECT 4.515 1.065 4.685 1.785 ;
        RECT 4.855 1.415 5.860 1.655 ;
        RECT 6.060 1.575 6.295 1.985 ;
        RECT 4.855 1.235 5.185 1.415 ;
        RECT 6.535 1.305 6.740 1.905 ;
        RECT 5.495 1.065 5.825 1.235 ;
        RECT 3.585 0.965 3.915 1.065 ;
        RECT 3.585 0.735 3.995 0.965 ;
        RECT 4.515 0.895 5.825 1.065 ;
        RECT 6.065 1.125 6.740 1.305 ;
        RECT 6.910 1.405 7.080 2.250 ;
        RECT 7.940 2.085 8.110 2.375 ;
        RECT 8.640 2.255 10.030 2.635 ;
        RECT 7.250 1.915 10.030 2.085 ;
        RECT 7.250 1.575 7.500 1.915 ;
        RECT 6.910 1.235 8.260 1.405 ;
        RECT 6.065 1.060 6.405 1.125 ;
        RECT 4.515 0.765 4.735 0.895 ;
        RECT 4.405 0.595 4.735 0.765 ;
        RECT 2.400 0.265 3.415 0.465 ;
        RECT 3.585 0.085 3.755 0.525 ;
        RECT 3.925 0.425 4.255 0.505 ;
        RECT 4.905 0.425 5.075 0.715 ;
        RECT 6.185 0.705 6.405 1.060 ;
        RECT 6.910 0.465 7.080 1.235 ;
        RECT 8.040 1.075 8.260 1.235 ;
        RECT 7.280 0.735 7.825 1.065 ;
        RECT 8.430 0.840 8.600 1.915 ;
        RECT 8.770 1.575 9.555 1.745 ;
        RECT 8.770 1.110 9.055 1.575 ;
        RECT 8.835 0.925 9.055 1.110 ;
        RECT 9.860 1.325 10.030 1.915 ;
        RECT 10.660 1.325 10.975 2.415 ;
        RECT 11.155 1.765 11.445 2.635 ;
        RECT 9.860 0.995 10.125 1.325 ;
        RECT 10.660 0.995 11.495 1.325 ;
        RECT 8.430 0.835 8.615 0.840 ;
        RECT 8.215 0.665 8.615 0.835 ;
        RECT 8.835 0.755 9.475 0.925 ;
        RECT 3.925 0.255 5.075 0.425 ;
        RECT 5.325 0.085 5.675 0.465 ;
        RECT 6.300 0.265 7.080 0.465 ;
        RECT 7.250 0.085 7.575 0.525 ;
        RECT 7.745 0.425 8.075 0.545 ;
        RECT 8.785 0.425 8.955 0.585 ;
        RECT 7.745 0.255 8.955 0.425 ;
        RECT 9.265 0.265 9.475 0.755 ;
        RECT 9.725 0.085 10.030 0.805 ;
        RECT 10.660 0.255 10.975 0.995 ;
        RECT 11.150 0.085 11.445 0.545 ;
        RECT 0.000 -0.085 11.960 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 0.610 0.765 0.780 0.935 ;
        RECT 1.065 1.785 1.235 1.955 ;
        RECT 2.445 1.785 2.615 1.955 ;
        RECT 2.905 0.765 3.075 0.935 ;
        RECT 6.125 1.785 6.295 1.955 ;
        RECT 5.665 1.445 5.835 1.615 ;
        RECT 3.825 0.765 3.995 0.935 ;
        RECT 6.125 1.105 6.295 1.275 ;
        RECT 7.575 0.765 7.745 0.935 ;
        RECT 8.855 1.445 9.025 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
      LAYER met1 ;
        RECT 1.005 1.940 1.295 1.985 ;
        RECT 2.385 1.940 2.675 1.985 ;
        RECT 6.065 1.940 6.355 1.985 ;
        RECT 1.005 1.800 6.355 1.940 ;
        RECT 1.005 1.755 1.295 1.800 ;
        RECT 2.385 1.755 2.675 1.800 ;
        RECT 6.065 1.755 6.355 1.800 ;
        RECT 5.605 1.600 5.895 1.645 ;
        RECT 8.795 1.600 9.085 1.645 ;
        RECT 5.605 1.460 9.085 1.600 ;
        RECT 5.605 1.415 5.895 1.460 ;
        RECT 8.795 1.415 9.085 1.460 ;
        RECT 6.065 1.260 6.355 1.305 ;
        RECT 2.920 1.120 6.355 1.260 ;
        RECT 2.920 0.965 3.135 1.120 ;
        RECT 6.065 1.075 6.355 1.120 ;
        RECT 0.550 0.920 0.840 0.965 ;
        RECT 2.845 0.920 3.135 0.965 ;
        RECT 0.550 0.780 3.135 0.920 ;
        RECT 0.550 0.735 0.840 0.780 ;
        RECT 2.845 0.735 3.135 0.780 ;
  END
END sky130_fd_sc_hd__dfbbn_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dfbbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfbbn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.440 1.625 ;
    END
  END CLK_N
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.760 1.005 2.170 1.625 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 9.250 1.095 9.730 1.325 ;
    END
  END RESET_B
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 3.780 0.920 4.070 0.965 ;
        RECT 7.460 0.920 7.750 0.965 ;
        RECT 3.780 0.780 7.750 0.920 ;
        RECT 3.780 0.735 4.070 0.780 ;
        RECT 7.460 0.735 7.750 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.880 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 9.650 1.005 12.875 1.015 ;
        RECT 3.920 0.785 6.190 1.005 ;
        RECT 7.795 0.785 12.875 1.005 ;
        RECT 0.005 0.105 12.875 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 13.070 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 12.880 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 12.115 1.445 12.345 2.465 ;
        RECT 12.160 0.825 12.345 1.445 ;
        RECT 12.115 0.255 12.345 0.825 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 10.240 1.630 10.500 2.465 ;
        RECT 10.320 0.715 10.500 1.630 ;
        RECT 10.240 0.255 10.500 0.715 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 12.880 2.805 ;
        RECT 0.085 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.085 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.085 0.635 0.840 0.805 ;
        RECT 0.085 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.240 2.465 ;
        RECT 1.445 2.135 1.785 2.635 ;
        RECT 1.955 1.965 2.125 2.465 ;
        RECT 2.350 2.250 3.180 2.420 ;
        RECT 1.420 1.795 2.125 1.965 ;
        RECT 1.420 0.825 1.590 1.795 ;
        RECT 2.340 1.575 2.840 1.955 ;
        RECT 1.420 0.635 2.125 0.825 ;
        RECT 2.340 0.705 2.560 1.575 ;
        RECT 3.010 1.405 3.180 2.250 ;
        RECT 3.420 2.205 3.800 2.635 ;
        RECT 4.100 2.035 4.270 2.375 ;
        RECT 3.350 1.785 4.700 2.035 ;
        RECT 4.890 1.915 5.220 2.635 ;
        RECT 6.265 2.250 7.095 2.420 ;
        RECT 7.335 2.255 7.715 2.635 ;
        RECT 3.350 1.575 3.600 1.785 ;
        RECT 4.110 1.405 4.360 1.485 ;
        RECT 3.010 1.235 4.360 1.405 ;
        RECT 3.010 1.195 3.410 1.235 ;
        RECT 2.740 0.645 3.070 1.015 ;
        RECT 1.445 0.085 1.785 0.465 ;
        RECT 1.955 0.305 2.125 0.635 ;
        RECT 3.240 0.465 3.410 1.195 ;
        RECT 4.140 1.155 4.360 1.235 ;
        RECT 4.530 1.065 4.700 1.785 ;
        RECT 4.870 1.415 5.875 1.655 ;
        RECT 6.075 1.575 6.310 1.985 ;
        RECT 4.870 1.235 5.200 1.415 ;
        RECT 6.550 1.305 6.755 1.905 ;
        RECT 5.510 1.065 5.840 1.235 ;
        RECT 3.600 0.965 3.930 1.065 ;
        RECT 3.600 0.735 4.010 0.965 ;
        RECT 4.530 0.895 5.840 1.065 ;
        RECT 6.135 1.125 6.755 1.305 ;
        RECT 6.925 1.405 7.095 2.250 ;
        RECT 7.955 2.085 8.125 2.375 ;
        RECT 8.655 2.255 10.070 2.635 ;
        RECT 7.265 1.915 10.070 2.085 ;
        RECT 7.265 1.575 7.515 1.915 ;
        RECT 6.925 1.235 8.275 1.405 ;
        RECT 4.530 0.765 4.750 0.895 ;
        RECT 4.420 0.595 4.750 0.765 ;
        RECT 2.415 0.265 3.410 0.465 ;
        RECT 3.580 0.085 3.750 0.525 ;
        RECT 3.920 0.425 4.250 0.545 ;
        RECT 4.920 0.425 5.170 0.715 ;
        RECT 6.135 0.705 6.420 1.125 ;
        RECT 6.925 0.465 7.095 1.235 ;
        RECT 8.055 1.075 8.275 1.235 ;
        RECT 7.470 0.735 7.845 1.065 ;
        RECT 8.445 0.780 8.625 1.915 ;
        RECT 8.295 0.595 8.625 0.780 ;
        RECT 8.795 1.575 9.570 1.745 ;
        RECT 8.795 0.925 9.070 1.575 ;
        RECT 9.900 1.325 10.070 1.915 ;
        RECT 10.680 1.465 10.910 2.635 ;
        RECT 11.215 1.325 11.470 2.415 ;
        RECT 11.650 1.765 11.945 2.635 ;
        RECT 12.515 1.465 12.795 2.635 ;
        RECT 9.900 0.995 10.140 1.325 ;
        RECT 11.215 0.995 11.990 1.325 ;
        RECT 8.795 0.755 9.500 0.925 ;
        RECT 3.920 0.255 5.170 0.425 ;
        RECT 5.360 0.085 5.690 0.465 ;
        RECT 6.330 0.265 7.095 0.465 ;
        RECT 7.275 0.085 7.535 0.525 ;
        RECT 7.795 0.425 8.125 0.545 ;
        RECT 8.795 0.425 8.965 0.585 ;
        RECT 7.795 0.255 8.965 0.425 ;
        RECT 9.280 0.265 9.500 0.755 ;
        RECT 9.740 0.085 10.070 0.805 ;
        RECT 10.680 0.085 10.910 0.885 ;
        RECT 11.215 0.255 11.470 0.995 ;
        RECT 11.650 0.085 11.945 0.545 ;
        RECT 12.515 0.085 12.795 0.885 ;
        RECT 0.000 -0.085 12.880 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 0.610 0.765 0.780 0.935 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.460 1.785 2.630 1.955 ;
        RECT 2.900 0.765 3.070 0.935 ;
        RECT 6.140 1.785 6.310 1.955 ;
        RECT 5.680 1.445 5.850 1.615 ;
        RECT 3.840 0.765 4.010 0.935 ;
        RECT 6.140 1.105 6.310 1.275 ;
        RECT 7.520 0.765 7.690 0.935 ;
        RECT 8.900 1.445 9.070 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.400 1.940 2.690 1.985 ;
        RECT 6.080 1.940 6.370 1.985 ;
        RECT 1.010 1.800 6.370 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.400 1.755 2.690 1.800 ;
        RECT 6.080 1.755 6.370 1.800 ;
        RECT 5.620 1.600 5.910 1.645 ;
        RECT 8.840 1.600 9.130 1.645 ;
        RECT 5.620 1.460 9.130 1.600 ;
        RECT 5.620 1.415 5.910 1.460 ;
        RECT 8.840 1.415 9.130 1.460 ;
        RECT 6.080 1.260 6.370 1.305 ;
        RECT 2.935 1.120 6.370 1.260 ;
        RECT 2.935 0.965 3.130 1.120 ;
        RECT 6.080 1.075 6.370 1.120 ;
        RECT 0.550 0.920 0.840 0.965 ;
        RECT 2.840 0.920 3.130 0.965 ;
        RECT 0.550 0.780 3.130 0.920 ;
        RECT 0.550 0.735 0.840 0.780 ;
        RECT 2.840 0.735 3.130 0.780 ;
  END
END sky130_fd_sc_hd__dfbbn_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dfbbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfbbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.960 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.750 1.005 2.160 1.625 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 9.315 1.095 9.690 1.325 ;
    END
  END RESET_B
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 3.770 0.920 4.060 0.965 ;
        RECT 7.450 0.920 7.740 0.965 ;
        RECT 3.770 0.780 7.740 0.920 ;
        RECT 3.770 0.735 4.060 0.780 ;
        RECT 7.450 0.735 7.740 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.960 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 9.620 1.005 11.955 1.015 ;
        RECT 3.910 0.785 6.180 1.005 ;
        RECT 7.785 0.785 11.955 1.005 ;
        RECT 0.005 0.105 11.955 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.150 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.960 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 11.615 1.445 11.875 2.465 ;
        RECT 11.660 0.825 11.875 1.445 ;
        RECT 11.615 0.255 11.875 0.825 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 10.200 1.630 10.485 2.465 ;
        RECT 10.280 0.715 10.485 1.630 ;
        RECT 10.200 0.255 10.485 0.715 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.960 2.805 ;
        RECT 0.085 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.085 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.085 0.635 0.840 0.805 ;
        RECT 0.085 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.240 2.465 ;
        RECT 1.435 2.135 1.785 2.635 ;
        RECT 1.955 1.965 2.125 2.465 ;
        RECT 2.340 2.250 3.170 2.420 ;
        RECT 1.410 1.795 2.125 1.965 ;
        RECT 1.410 0.825 1.580 1.795 ;
        RECT 2.330 1.575 2.830 1.955 ;
        RECT 1.410 0.635 2.125 0.825 ;
        RECT 2.330 0.705 2.550 1.575 ;
        RECT 3.000 1.405 3.170 2.250 ;
        RECT 3.410 2.205 3.790 2.635 ;
        RECT 4.090 2.035 4.260 2.375 ;
        RECT 3.340 1.785 4.690 2.035 ;
        RECT 4.880 1.915 5.210 2.635 ;
        RECT 6.255 2.250 7.085 2.420 ;
        RECT 7.325 2.255 7.705 2.635 ;
        RECT 3.340 1.575 3.590 1.785 ;
        RECT 4.100 1.405 4.350 1.485 ;
        RECT 3.000 1.235 4.350 1.405 ;
        RECT 3.000 1.195 3.400 1.235 ;
        RECT 2.730 0.645 3.060 1.015 ;
        RECT 1.435 0.085 1.785 0.465 ;
        RECT 1.955 0.305 2.125 0.635 ;
        RECT 3.230 0.465 3.400 1.195 ;
        RECT 4.130 1.155 4.350 1.235 ;
        RECT 4.520 1.065 4.690 1.785 ;
        RECT 4.860 1.415 5.865 1.655 ;
        RECT 6.065 1.575 6.300 1.985 ;
        RECT 4.860 1.235 5.190 1.415 ;
        RECT 6.540 1.305 6.745 1.905 ;
        RECT 5.500 1.065 5.830 1.235 ;
        RECT 3.590 0.965 3.920 1.065 ;
        RECT 3.590 0.735 4.000 0.965 ;
        RECT 4.520 0.895 5.830 1.065 ;
        RECT 6.125 1.125 6.745 1.305 ;
        RECT 6.915 1.405 7.085 2.250 ;
        RECT 7.945 2.085 8.115 2.375 ;
        RECT 8.645 2.255 10.030 2.635 ;
        RECT 7.255 1.915 10.030 2.085 ;
        RECT 7.255 1.575 7.505 1.915 ;
        RECT 6.915 1.235 8.265 1.405 ;
        RECT 4.520 0.765 4.740 0.895 ;
        RECT 4.410 0.595 4.740 0.765 ;
        RECT 2.405 0.265 3.400 0.465 ;
        RECT 3.570 0.085 3.740 0.525 ;
        RECT 3.910 0.425 4.240 0.545 ;
        RECT 4.910 0.425 5.080 0.715 ;
        RECT 6.125 0.705 6.410 1.125 ;
        RECT 6.915 0.465 7.085 1.235 ;
        RECT 8.045 1.075 8.265 1.235 ;
        RECT 7.460 0.735 7.835 1.065 ;
        RECT 8.435 0.780 8.615 1.915 ;
        RECT 8.285 0.595 8.615 0.780 ;
        RECT 8.785 1.575 9.545 1.745 ;
        RECT 8.785 0.925 9.060 1.575 ;
        RECT 9.860 1.325 10.030 1.915 ;
        RECT 10.655 1.325 10.970 2.415 ;
        RECT 11.150 1.765 11.445 2.635 ;
        RECT 9.860 0.995 10.110 1.325 ;
        RECT 10.655 0.995 11.490 1.325 ;
        RECT 8.785 0.755 9.475 0.925 ;
        RECT 3.910 0.255 5.080 0.425 ;
        RECT 5.350 0.085 5.680 0.465 ;
        RECT 6.320 0.265 7.085 0.465 ;
        RECT 7.265 0.085 7.525 0.525 ;
        RECT 7.785 0.425 8.115 0.545 ;
        RECT 8.785 0.425 8.955 0.585 ;
        RECT 7.785 0.255 8.955 0.425 ;
        RECT 9.240 0.265 9.475 0.755 ;
        RECT 9.700 0.085 10.030 0.805 ;
        RECT 10.655 0.255 10.970 0.995 ;
        RECT 11.150 0.085 11.445 0.545 ;
        RECT 0.000 -0.085 11.960 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 0.610 1.785 0.780 1.955 ;
        RECT 1.070 0.765 1.240 0.935 ;
        RECT 2.450 1.785 2.620 1.955 ;
        RECT 2.890 0.765 3.060 0.935 ;
        RECT 6.130 1.785 6.300 1.955 ;
        RECT 5.670 1.445 5.840 1.615 ;
        RECT 3.830 0.765 4.000 0.935 ;
        RECT 6.130 1.105 6.300 1.275 ;
        RECT 7.510 0.765 7.680 0.935 ;
        RECT 8.890 1.445 9.060 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
      LAYER met1 ;
        RECT 0.550 1.940 0.840 1.985 ;
        RECT 2.390 1.940 2.680 1.985 ;
        RECT 6.070 1.940 6.360 1.985 ;
        RECT 0.550 1.800 6.360 1.940 ;
        RECT 0.550 1.755 0.840 1.800 ;
        RECT 2.390 1.755 2.680 1.800 ;
        RECT 6.070 1.755 6.360 1.800 ;
        RECT 5.610 1.600 5.900 1.645 ;
        RECT 8.830 1.600 9.120 1.645 ;
        RECT 5.610 1.460 9.120 1.600 ;
        RECT 5.610 1.415 5.900 1.460 ;
        RECT 8.830 1.415 9.120 1.460 ;
        RECT 6.070 1.260 6.360 1.305 ;
        RECT 2.925 1.120 6.360 1.260 ;
        RECT 2.925 0.965 3.120 1.120 ;
        RECT 6.070 1.075 6.360 1.120 ;
        RECT 1.010 0.920 1.300 0.965 ;
        RECT 2.830 0.920 3.120 0.965 ;
        RECT 1.010 0.780 3.120 0.920 ;
        RECT 1.010 0.735 1.300 0.780 ;
        RECT 2.830 0.735 3.120 0.780 ;
  END
END sky130_fd_sc_hd__dfbbp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.580 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.680 2.450 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 7.045 0.965 7.335 1.280 ;
        RECT 3.745 0.920 4.395 0.965 ;
        RECT 7.045 0.920 7.635 0.965 ;
        RECT 3.745 0.780 7.635 0.920 ;
        RECT 3.745 0.735 4.395 0.780 ;
        RECT 7.345 0.735 7.635 0.780 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.580 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.515 0.785 5.445 1.005 ;
        RECT 8.165 0.785 10.520 1.015 ;
        RECT 0.005 0.105 10.520 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.770 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.580 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.449000 ;
    PORT
      LAYER li1 ;
        RECT 8.600 1.455 9.005 2.465 ;
        RECT 8.675 0.275 9.005 1.455 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 10.180 1.445 10.435 2.325 ;
        RECT 10.225 0.795 10.435 1.445 ;
        RECT 10.180 0.265 10.435 0.795 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.580 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.090 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.090 0.635 0.840 0.805 ;
        RECT 0.090 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 2.465 ;
        RECT 1.850 2.175 2.100 2.635 ;
        RECT 2.270 2.135 2.520 2.465 ;
        RECT 2.735 2.135 3.415 2.465 ;
        RECT 2.270 2.005 2.440 2.135 ;
        RECT 2.045 1.835 2.440 2.005 ;
        RECT 2.045 0.475 2.215 1.835 ;
        RECT 2.610 1.575 3.075 1.965 ;
        RECT 2.385 0.765 2.735 1.385 ;
        RECT 2.905 0.985 3.075 1.575 ;
        RECT 3.245 1.355 3.415 2.135 ;
        RECT 3.585 2.035 3.755 2.375 ;
        RECT 3.990 2.205 4.320 2.635 ;
        RECT 4.490 2.035 4.660 2.375 ;
        RECT 4.955 2.175 5.325 2.635 ;
        RECT 3.585 1.865 4.660 2.035 ;
        RECT 5.495 2.005 5.665 2.465 ;
        RECT 5.900 2.125 6.770 2.465 ;
        RECT 6.940 2.175 7.190 2.635 ;
        RECT 5.105 1.835 5.665 2.005 ;
        RECT 5.105 1.695 5.275 1.835 ;
        RECT 3.775 1.525 5.275 1.695 ;
        RECT 5.970 1.665 6.430 1.955 ;
        RECT 3.245 1.185 4.935 1.355 ;
        RECT 2.905 0.765 3.260 0.985 ;
        RECT 3.430 0.475 3.600 1.185 ;
        RECT 3.805 0.765 4.595 1.015 ;
        RECT 4.765 1.005 4.935 1.185 ;
        RECT 5.105 0.835 5.275 1.525 ;
        RECT 1.545 0.085 1.875 0.445 ;
        RECT 2.045 0.305 2.540 0.475 ;
        RECT 2.745 0.305 3.600 0.475 ;
        RECT 4.475 0.085 4.805 0.545 ;
        RECT 5.015 0.445 5.275 0.835 ;
        RECT 5.465 1.655 6.430 1.665 ;
        RECT 6.600 1.745 6.770 2.125 ;
        RECT 7.360 2.085 7.530 2.375 ;
        RECT 7.710 2.255 8.430 2.635 ;
        RECT 7.360 1.915 8.160 2.085 ;
        RECT 5.465 1.495 6.140 1.655 ;
        RECT 6.600 1.575 7.820 1.745 ;
        RECT 5.465 0.705 5.675 1.495 ;
        RECT 6.600 1.485 6.770 1.575 ;
        RECT 5.845 0.705 6.195 1.325 ;
        RECT 6.365 1.315 6.770 1.485 ;
        RECT 6.365 0.535 6.535 1.315 ;
        RECT 6.705 0.865 6.925 1.145 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.990 1.325 8.160 1.915 ;
        RECT 9.195 1.325 9.525 2.425 ;
        RECT 9.760 1.495 9.930 2.635 ;
        RECT 7.990 1.295 8.435 1.325 ;
        RECT 6.705 0.695 7.235 0.865 ;
        RECT 5.015 0.275 5.365 0.445 ;
        RECT 5.585 0.255 6.535 0.535 ;
        RECT 6.705 0.085 6.895 0.525 ;
        RECT 7.065 0.465 7.235 0.695 ;
        RECT 7.405 0.635 7.645 1.035 ;
        RECT 7.815 0.995 8.435 1.295 ;
        RECT 9.195 0.995 10.055 1.325 ;
        RECT 7.815 0.820 8.140 0.995 ;
        RECT 7.815 0.465 8.135 0.820 ;
        RECT 7.065 0.295 8.135 0.465 ;
        RECT 8.335 0.085 8.505 0.770 ;
        RECT 9.195 0.345 9.445 0.995 ;
        RECT 9.760 0.085 9.930 0.680 ;
        RECT 0.000 -0.085 10.580 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 0.610 1.105 0.780 1.275 ;
        RECT 1.015 1.785 1.185 1.955 ;
        RECT 2.905 1.785 3.075 1.955 ;
        RECT 2.445 1.105 2.615 1.275 ;
        RECT 6.025 1.785 6.195 1.955 ;
        RECT 4.165 0.765 4.335 0.935 ;
        RECT 6.025 1.105 6.195 1.275 ;
        RECT 7.105 1.080 7.275 1.250 ;
        RECT 7.405 0.765 7.575 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
      LAYER met1 ;
        RECT 0.955 1.940 1.245 1.985 ;
        RECT 2.845 1.940 3.135 1.985 ;
        RECT 5.965 1.940 6.255 1.985 ;
        RECT 0.955 1.800 6.255 1.940 ;
        RECT 0.955 1.755 1.245 1.800 ;
        RECT 2.845 1.755 3.135 1.800 ;
        RECT 5.965 1.755 6.255 1.800 ;
        RECT 0.550 1.260 0.840 1.305 ;
        RECT 2.385 1.260 2.675 1.305 ;
        RECT 5.965 1.260 6.255 1.305 ;
        RECT 0.550 1.120 6.255 1.260 ;
        RECT 0.550 1.075 0.840 1.120 ;
        RECT 2.385 1.075 2.675 1.120 ;
        RECT 5.965 1.075 6.255 1.120 ;
  END
END sky130_fd_sc_hd__dfrbp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dfrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.680 2.450 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 7.045 0.965 7.335 1.280 ;
        RECT 3.745 0.920 4.395 0.965 ;
        RECT 7.045 0.920 7.635 0.965 ;
        RECT 3.745 0.780 7.635 0.920 ;
        RECT 3.745 0.735 4.395 0.780 ;
        RECT 7.345 0.735 7.635 0.780 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.515 0.785 5.445 1.005 ;
        RECT 8.650 0.785 10.930 1.015 ;
        RECT 0.005 0.105 10.930 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.511500 ;
    PORT
      LAYER li1 ;
        RECT 9.160 0.265 9.495 1.695 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 10.120 2.080 10.420 2.465 ;
        RECT 10.030 1.535 10.420 2.080 ;
        RECT 10.250 0.825 10.420 1.535 ;
        RECT 10.040 0.310 10.420 0.825 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.090 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.090 0.635 0.840 0.805 ;
        RECT 0.090 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 2.465 ;
        RECT 1.850 2.175 2.100 2.635 ;
        RECT 2.270 2.135 2.520 2.465 ;
        RECT 2.735 2.135 3.415 2.465 ;
        RECT 2.270 2.005 2.440 2.135 ;
        RECT 2.045 1.835 2.440 2.005 ;
        RECT 2.045 0.475 2.215 1.835 ;
        RECT 2.610 1.575 3.075 1.965 ;
        RECT 2.385 0.765 2.735 1.385 ;
        RECT 2.905 0.985 3.075 1.575 ;
        RECT 3.245 1.355 3.415 2.135 ;
        RECT 3.585 2.035 3.755 2.375 ;
        RECT 3.990 2.205 4.320 2.635 ;
        RECT 4.490 2.035 4.660 2.375 ;
        RECT 4.955 2.175 5.325 2.635 ;
        RECT 3.585 1.865 4.660 2.035 ;
        RECT 5.495 2.005 5.665 2.465 ;
        RECT 5.900 2.125 6.770 2.465 ;
        RECT 6.940 2.175 7.190 2.635 ;
        RECT 5.105 1.835 5.665 2.005 ;
        RECT 5.105 1.695 5.275 1.835 ;
        RECT 3.775 1.525 5.275 1.695 ;
        RECT 5.970 1.665 6.430 1.955 ;
        RECT 3.245 1.185 4.935 1.355 ;
        RECT 2.905 0.765 3.260 0.985 ;
        RECT 3.430 0.475 3.600 1.185 ;
        RECT 3.805 0.765 4.595 1.015 ;
        RECT 4.765 1.005 4.935 1.185 ;
        RECT 5.105 0.835 5.275 1.525 ;
        RECT 1.545 0.085 1.875 0.445 ;
        RECT 2.045 0.305 2.540 0.475 ;
        RECT 2.745 0.305 3.600 0.475 ;
        RECT 4.475 0.085 4.805 0.545 ;
        RECT 5.015 0.445 5.275 0.835 ;
        RECT 5.465 1.655 6.430 1.665 ;
        RECT 6.600 1.745 6.770 2.125 ;
        RECT 7.360 2.085 7.530 2.375 ;
        RECT 7.710 2.255 8.055 2.635 ;
        RECT 7.360 1.915 8.160 2.085 ;
        RECT 5.465 1.495 6.140 1.655 ;
        RECT 6.600 1.575 7.820 1.745 ;
        RECT 5.465 0.705 5.675 1.495 ;
        RECT 6.600 1.485 6.770 1.575 ;
        RECT 5.845 0.705 6.195 1.325 ;
        RECT 6.365 1.315 6.770 1.485 ;
        RECT 6.365 0.535 6.535 1.315 ;
        RECT 6.705 0.865 6.925 1.145 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.990 1.325 8.160 1.915 ;
        RECT 8.335 2.035 8.560 2.465 ;
        RECT 8.730 2.205 9.070 2.635 ;
        RECT 9.620 2.255 9.950 2.635 ;
        RECT 8.335 1.865 9.835 2.035 ;
        RECT 8.335 1.795 8.990 1.865 ;
        RECT 7.990 1.295 8.650 1.325 ;
        RECT 6.705 0.695 7.235 0.865 ;
        RECT 5.015 0.275 5.365 0.445 ;
        RECT 5.585 0.255 6.535 0.535 ;
        RECT 6.705 0.085 6.895 0.525 ;
        RECT 7.065 0.465 7.235 0.695 ;
        RECT 7.405 0.635 7.645 1.035 ;
        RECT 7.815 1.075 8.650 1.295 ;
        RECT 7.815 0.995 8.160 1.075 ;
        RECT 7.815 0.465 7.985 0.995 ;
        RECT 8.820 0.885 8.990 1.795 ;
        RECT 9.665 1.325 9.835 1.865 ;
        RECT 10.590 1.445 10.760 2.635 ;
        RECT 9.665 0.995 10.080 1.325 ;
        RECT 7.065 0.295 7.985 0.465 ;
        RECT 8.335 0.715 8.990 0.885 ;
        RECT 8.335 0.345 8.585 0.715 ;
        RECT 8.755 0.085 8.990 0.545 ;
        RECT 9.700 0.085 9.870 0.825 ;
        RECT 10.590 0.085 10.760 0.930 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 0.610 1.105 0.780 1.275 ;
        RECT 1.015 1.785 1.185 1.955 ;
        RECT 2.905 1.785 3.075 1.955 ;
        RECT 2.445 1.105 2.615 1.275 ;
        RECT 6.025 1.785 6.195 1.955 ;
        RECT 4.165 0.765 4.335 0.935 ;
        RECT 6.025 1.105 6.195 1.275 ;
        RECT 7.105 1.080 7.275 1.250 ;
        RECT 7.405 0.765 7.575 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
      LAYER met1 ;
        RECT 0.955 1.940 1.245 1.985 ;
        RECT 2.845 1.940 3.135 1.985 ;
        RECT 5.965 1.940 6.255 1.985 ;
        RECT 0.955 1.800 6.255 1.940 ;
        RECT 0.955 1.755 1.245 1.800 ;
        RECT 2.845 1.755 3.135 1.800 ;
        RECT 5.965 1.755 6.255 1.800 ;
        RECT 0.550 1.260 0.840 1.305 ;
        RECT 2.385 1.260 2.675 1.305 ;
        RECT 5.965 1.260 6.255 1.305 ;
        RECT 0.550 1.120 6.255 1.260 ;
        RECT 0.550 1.075 0.840 1.120 ;
        RECT 2.385 1.075 2.675 1.120 ;
        RECT 5.965 1.075 6.255 1.120 ;
  END
END sky130_fd_sc_hd__dfrbp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dfrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK_N
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.680 2.450 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 7.045 0.965 7.335 1.280 ;
        RECT 3.745 0.920 4.395 0.965 ;
        RECT 7.045 0.920 7.635 0.965 ;
        RECT 3.745 0.780 7.635 0.920 ;
        RECT 3.745 0.735 4.395 0.780 ;
        RECT 7.345 0.735 7.635 0.780 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.515 0.785 5.445 1.005 ;
        RECT 8.275 0.785 9.195 1.015 ;
        RECT 0.005 0.105 9.195 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.390 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 8.855 1.445 9.110 2.325 ;
        RECT 8.900 0.795 9.110 1.445 ;
        RECT 8.855 0.265 9.110 0.795 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.090 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.090 0.635 0.840 0.805 ;
        RECT 0.090 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 2.465 ;
        RECT 1.850 2.175 2.100 2.635 ;
        RECT 2.270 2.135 2.520 2.465 ;
        RECT 2.735 2.135 3.415 2.465 ;
        RECT 2.270 2.005 2.440 2.135 ;
        RECT 2.045 1.835 2.440 2.005 ;
        RECT 2.045 0.475 2.215 1.835 ;
        RECT 2.610 1.575 3.075 1.965 ;
        RECT 2.385 0.765 2.735 1.385 ;
        RECT 2.905 0.985 3.075 1.575 ;
        RECT 3.245 1.355 3.415 2.135 ;
        RECT 3.585 2.035 3.755 2.375 ;
        RECT 3.990 2.205 4.320 2.635 ;
        RECT 4.490 2.035 4.660 2.375 ;
        RECT 4.955 2.175 5.325 2.635 ;
        RECT 3.585 1.865 4.660 2.035 ;
        RECT 5.495 2.005 5.665 2.465 ;
        RECT 5.900 2.125 6.770 2.465 ;
        RECT 6.940 2.175 7.190 2.635 ;
        RECT 5.105 1.835 5.665 2.005 ;
        RECT 5.105 1.695 5.275 1.835 ;
        RECT 3.775 1.525 5.275 1.695 ;
        RECT 5.970 1.665 6.430 1.955 ;
        RECT 3.245 1.185 4.935 1.355 ;
        RECT 2.905 0.765 3.260 0.985 ;
        RECT 3.430 0.475 3.600 1.185 ;
        RECT 3.805 0.765 4.595 1.015 ;
        RECT 4.765 1.005 4.935 1.185 ;
        RECT 5.105 0.835 5.275 1.525 ;
        RECT 1.545 0.085 1.875 0.445 ;
        RECT 2.045 0.305 2.540 0.475 ;
        RECT 2.745 0.305 3.600 0.475 ;
        RECT 4.475 0.085 4.805 0.545 ;
        RECT 5.015 0.445 5.275 0.835 ;
        RECT 5.465 1.655 6.430 1.665 ;
        RECT 6.600 1.745 6.770 2.125 ;
        RECT 7.360 2.085 7.530 2.375 ;
        RECT 7.710 2.255 8.040 2.635 ;
        RECT 7.360 1.915 8.160 2.085 ;
        RECT 5.465 1.495 6.140 1.655 ;
        RECT 6.600 1.575 7.820 1.745 ;
        RECT 5.465 0.705 5.675 1.495 ;
        RECT 6.600 1.485 6.770 1.575 ;
        RECT 5.845 0.705 6.195 1.325 ;
        RECT 6.365 1.315 6.770 1.485 ;
        RECT 6.365 0.535 6.535 1.315 ;
        RECT 6.705 0.865 6.925 1.145 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.990 1.325 8.160 1.915 ;
        RECT 8.380 1.495 8.685 2.635 ;
        RECT 7.990 1.295 8.730 1.325 ;
        RECT 6.705 0.695 7.235 0.865 ;
        RECT 5.015 0.275 5.365 0.445 ;
        RECT 5.585 0.255 6.535 0.535 ;
        RECT 6.705 0.085 6.895 0.525 ;
        RECT 7.065 0.465 7.235 0.695 ;
        RECT 7.405 0.635 7.645 1.035 ;
        RECT 7.815 0.995 8.730 1.295 ;
        RECT 7.815 0.820 8.140 0.995 ;
        RECT 7.815 0.465 8.135 0.820 ;
        RECT 7.065 0.295 8.135 0.465 ;
        RECT 8.380 0.085 8.685 0.545 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 0.655 1.785 0.825 1.955 ;
        RECT 1.015 1.105 1.185 1.275 ;
        RECT 2.905 1.785 3.075 1.955 ;
        RECT 2.445 1.105 2.615 1.275 ;
        RECT 6.025 1.785 6.195 1.955 ;
        RECT 4.165 0.765 4.335 0.935 ;
        RECT 6.025 1.105 6.195 1.275 ;
        RECT 7.105 1.080 7.275 1.250 ;
        RECT 7.405 0.765 7.575 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
      LAYER met1 ;
        RECT 0.595 1.940 0.885 1.985 ;
        RECT 2.845 1.940 3.135 1.985 ;
        RECT 5.965 1.940 6.255 1.985 ;
        RECT 0.595 1.800 6.255 1.940 ;
        RECT 0.595 1.755 0.885 1.800 ;
        RECT 2.845 1.755 3.135 1.800 ;
        RECT 5.965 1.755 6.255 1.800 ;
        RECT 0.955 1.260 1.245 1.305 ;
        RECT 2.385 1.260 2.675 1.305 ;
        RECT 5.965 1.260 6.255 1.305 ;
        RECT 0.955 1.120 6.255 1.260 ;
        RECT 0.955 1.075 1.245 1.120 ;
        RECT 2.385 1.075 2.675 1.120 ;
        RECT 5.965 1.075 6.255 1.120 ;
  END
END sky130_fd_sc_hd__dfrtn_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.680 2.450 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 7.045 0.965 7.335 1.280 ;
        RECT 3.745 0.920 4.395 0.965 ;
        RECT 7.045 0.920 7.635 0.965 ;
        RECT 3.745 0.780 7.635 0.920 ;
        RECT 3.745 0.735 4.395 0.780 ;
        RECT 7.345 0.735 7.635 0.780 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.515 0.785 5.445 1.005 ;
        RECT 8.275 0.785 9.195 1.015 ;
        RECT 0.005 0.105 9.195 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.390 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 8.855 1.445 9.110 2.325 ;
        RECT 8.900 0.795 9.110 1.445 ;
        RECT 8.855 0.265 9.110 0.795 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.090 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.090 0.635 0.840 0.805 ;
        RECT 0.090 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 2.465 ;
        RECT 1.850 2.175 2.100 2.635 ;
        RECT 2.270 2.135 2.520 2.465 ;
        RECT 2.735 2.135 3.415 2.465 ;
        RECT 2.270 2.005 2.440 2.135 ;
        RECT 2.045 1.835 2.440 2.005 ;
        RECT 2.045 0.475 2.215 1.835 ;
        RECT 2.610 1.575 3.075 1.965 ;
        RECT 2.385 0.765 2.735 1.385 ;
        RECT 2.905 0.985 3.075 1.575 ;
        RECT 3.245 1.355 3.415 2.135 ;
        RECT 3.585 2.035 3.755 2.375 ;
        RECT 3.990 2.205 4.320 2.635 ;
        RECT 4.490 2.035 4.660 2.375 ;
        RECT 4.955 2.175 5.325 2.635 ;
        RECT 3.585 1.865 4.660 2.035 ;
        RECT 5.495 2.005 5.665 2.465 ;
        RECT 5.900 2.125 6.770 2.465 ;
        RECT 6.940 2.175 7.190 2.635 ;
        RECT 5.105 1.835 5.665 2.005 ;
        RECT 5.105 1.695 5.275 1.835 ;
        RECT 3.775 1.525 5.275 1.695 ;
        RECT 5.970 1.665 6.430 1.955 ;
        RECT 3.245 1.185 4.935 1.355 ;
        RECT 2.905 0.765 3.260 0.985 ;
        RECT 3.430 0.475 3.600 1.185 ;
        RECT 3.805 0.765 4.595 1.015 ;
        RECT 4.765 1.005 4.935 1.185 ;
        RECT 5.105 0.835 5.275 1.525 ;
        RECT 1.545 0.085 1.875 0.445 ;
        RECT 2.045 0.305 2.540 0.475 ;
        RECT 2.745 0.305 3.600 0.475 ;
        RECT 4.475 0.085 4.805 0.545 ;
        RECT 5.015 0.445 5.275 0.835 ;
        RECT 5.465 1.655 6.430 1.665 ;
        RECT 6.600 1.745 6.770 2.125 ;
        RECT 7.360 2.085 7.530 2.375 ;
        RECT 7.710 2.255 8.040 2.635 ;
        RECT 7.360 1.915 8.160 2.085 ;
        RECT 5.465 1.495 6.140 1.655 ;
        RECT 6.600 1.575 7.820 1.745 ;
        RECT 5.465 0.705 5.675 1.495 ;
        RECT 6.600 1.485 6.770 1.575 ;
        RECT 5.845 0.705 6.195 1.325 ;
        RECT 6.365 1.315 6.770 1.485 ;
        RECT 6.365 0.535 6.535 1.315 ;
        RECT 6.705 0.865 6.925 1.145 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.990 1.325 8.160 1.915 ;
        RECT 8.380 1.495 8.685 2.635 ;
        RECT 7.990 1.295 8.730 1.325 ;
        RECT 6.705 0.695 7.235 0.865 ;
        RECT 5.015 0.275 5.365 0.445 ;
        RECT 5.585 0.255 6.535 0.535 ;
        RECT 6.705 0.085 6.895 0.525 ;
        RECT 7.065 0.465 7.235 0.695 ;
        RECT 7.405 0.635 7.645 1.035 ;
        RECT 7.815 0.995 8.730 1.295 ;
        RECT 7.815 0.820 8.140 0.995 ;
        RECT 7.815 0.465 8.135 0.820 ;
        RECT 7.065 0.295 8.135 0.465 ;
        RECT 8.380 0.085 8.685 0.545 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 0.610 1.105 0.780 1.275 ;
        RECT 1.015 1.785 1.185 1.955 ;
        RECT 2.905 1.785 3.075 1.955 ;
        RECT 2.445 1.105 2.615 1.275 ;
        RECT 6.025 1.785 6.195 1.955 ;
        RECT 4.165 0.765 4.335 0.935 ;
        RECT 6.025 1.105 6.195 1.275 ;
        RECT 7.105 1.080 7.275 1.250 ;
        RECT 7.405 0.765 7.575 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
      LAYER met1 ;
        RECT 0.955 1.940 1.245 1.985 ;
        RECT 2.845 1.940 3.135 1.985 ;
        RECT 5.965 1.940 6.255 1.985 ;
        RECT 0.955 1.800 6.255 1.940 ;
        RECT 0.955 1.755 1.245 1.800 ;
        RECT 2.845 1.755 3.135 1.800 ;
        RECT 5.965 1.755 6.255 1.800 ;
        RECT 0.550 1.260 0.840 1.305 ;
        RECT 2.385 1.260 2.675 1.305 ;
        RECT 5.965 1.260 6.255 1.305 ;
        RECT 0.550 1.120 6.255 1.260 ;
        RECT 0.550 1.075 0.840 1.120 ;
        RECT 2.385 1.075 2.675 1.120 ;
        RECT 5.965 1.075 6.255 1.120 ;
  END
END sky130_fd_sc_hd__dfrtp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dfrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.680 2.450 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 7.045 0.965 7.335 1.280 ;
        RECT 3.745 0.920 4.395 0.965 ;
        RECT 7.045 0.920 7.635 0.965 ;
        RECT 3.745 0.780 7.635 0.920 ;
        RECT 3.745 0.735 4.395 0.780 ;
        RECT 7.345 0.735 7.635 0.780 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.515 0.785 5.445 1.005 ;
        RECT 8.275 0.785 9.615 1.015 ;
        RECT 0.005 0.105 9.615 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 8.855 1.445 9.105 2.325 ;
        RECT 8.900 0.795 9.105 1.445 ;
        RECT 8.855 0.265 9.105 0.795 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.090 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.090 0.635 0.840 0.805 ;
        RECT 0.090 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 2.465 ;
        RECT 1.850 2.175 2.100 2.635 ;
        RECT 2.270 2.135 2.520 2.465 ;
        RECT 2.735 2.135 3.415 2.465 ;
        RECT 2.270 2.005 2.440 2.135 ;
        RECT 2.045 1.835 2.440 2.005 ;
        RECT 2.045 0.475 2.215 1.835 ;
        RECT 2.610 1.575 3.075 1.965 ;
        RECT 2.385 0.765 2.735 1.385 ;
        RECT 2.905 0.985 3.075 1.575 ;
        RECT 3.245 1.355 3.415 2.135 ;
        RECT 3.585 2.035 3.755 2.375 ;
        RECT 3.990 2.205 4.320 2.635 ;
        RECT 4.490 2.035 4.660 2.375 ;
        RECT 4.955 2.175 5.325 2.635 ;
        RECT 3.585 1.865 4.660 2.035 ;
        RECT 5.495 2.005 5.665 2.465 ;
        RECT 5.900 2.125 6.770 2.465 ;
        RECT 6.940 2.175 7.190 2.635 ;
        RECT 5.105 1.835 5.665 2.005 ;
        RECT 5.105 1.695 5.275 1.835 ;
        RECT 3.775 1.525 5.275 1.695 ;
        RECT 5.970 1.665 6.430 1.955 ;
        RECT 3.245 1.185 4.935 1.355 ;
        RECT 2.905 0.765 3.260 0.985 ;
        RECT 3.430 0.475 3.600 1.185 ;
        RECT 3.805 0.765 4.595 1.015 ;
        RECT 4.765 1.005 4.935 1.185 ;
        RECT 5.105 0.835 5.275 1.525 ;
        RECT 1.545 0.085 1.875 0.445 ;
        RECT 2.045 0.305 2.540 0.475 ;
        RECT 2.745 0.305 3.600 0.475 ;
        RECT 4.475 0.085 4.805 0.545 ;
        RECT 5.015 0.445 5.275 0.835 ;
        RECT 5.465 1.655 6.430 1.665 ;
        RECT 6.600 1.745 6.770 2.125 ;
        RECT 7.360 2.085 7.530 2.375 ;
        RECT 7.710 2.255 8.040 2.635 ;
        RECT 7.360 1.915 8.160 2.085 ;
        RECT 5.465 1.495 6.140 1.655 ;
        RECT 6.600 1.575 7.820 1.745 ;
        RECT 5.465 0.705 5.675 1.495 ;
        RECT 6.600 1.485 6.770 1.575 ;
        RECT 5.845 0.705 6.195 1.325 ;
        RECT 6.365 1.315 6.770 1.485 ;
        RECT 6.365 0.535 6.535 1.315 ;
        RECT 6.705 0.865 6.925 1.145 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.990 1.325 8.160 1.915 ;
        RECT 8.380 1.495 8.685 2.635 ;
        RECT 9.275 1.495 9.525 2.635 ;
        RECT 7.990 1.295 8.730 1.325 ;
        RECT 6.705 0.695 7.235 0.865 ;
        RECT 5.015 0.275 5.365 0.445 ;
        RECT 5.585 0.255 6.535 0.535 ;
        RECT 6.705 0.085 6.895 0.525 ;
        RECT 7.065 0.465 7.235 0.695 ;
        RECT 7.405 0.635 7.645 1.035 ;
        RECT 7.815 0.995 8.730 1.295 ;
        RECT 7.815 0.820 8.140 0.995 ;
        RECT 7.815 0.465 8.135 0.820 ;
        RECT 7.065 0.295 8.135 0.465 ;
        RECT 8.380 0.085 8.685 0.545 ;
        RECT 9.275 0.085 9.525 0.840 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.610 1.105 0.780 1.275 ;
        RECT 1.015 1.785 1.185 1.955 ;
        RECT 2.905 1.785 3.075 1.955 ;
        RECT 2.445 1.105 2.615 1.275 ;
        RECT 6.025 1.785 6.195 1.955 ;
        RECT 4.165 0.765 4.335 0.935 ;
        RECT 6.025 1.105 6.195 1.275 ;
        RECT 7.105 1.080 7.275 1.250 ;
        RECT 7.405 0.765 7.575 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 0.955 1.940 1.245 1.985 ;
        RECT 2.845 1.940 3.135 1.985 ;
        RECT 5.965 1.940 6.255 1.985 ;
        RECT 0.955 1.800 6.255 1.940 ;
        RECT 0.955 1.755 1.245 1.800 ;
        RECT 2.845 1.755 3.135 1.800 ;
        RECT 5.965 1.755 6.255 1.800 ;
        RECT 0.550 1.260 0.840 1.305 ;
        RECT 2.385 1.260 2.675 1.305 ;
        RECT 5.965 1.260 6.255 1.305 ;
        RECT 0.550 1.120 6.255 1.260 ;
        RECT 0.550 1.075 0.840 1.120 ;
        RECT 2.385 1.075 2.675 1.120 ;
        RECT 5.965 1.075 6.255 1.120 ;
  END
END sky130_fd_sc_hd__dfrtp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dfrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfrtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.580 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.355 1.665 1.680 2.450 ;
        RECT 1.415 0.615 1.875 1.665 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 7.045 0.965 7.335 1.280 ;
        RECT 3.745 0.920 4.395 0.965 ;
        RECT 7.045 0.920 7.635 0.965 ;
        RECT 3.745 0.780 7.635 0.920 ;
        RECT 3.745 0.735 4.395 0.780 ;
        RECT 7.345 0.735 7.635 0.780 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.580 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.515 0.785 5.445 1.005 ;
        RECT 8.165 0.785 10.375 1.015 ;
        RECT 0.005 0.105 10.375 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.770 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.580 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 8.715 1.625 9.005 2.465 ;
        RECT 9.555 1.625 9.805 2.465 ;
        RECT 8.715 1.455 10.440 1.625 ;
        RECT 10.030 0.905 10.440 1.455 ;
        RECT 8.675 0.735 10.440 0.905 ;
        RECT 8.675 0.255 9.005 0.735 ;
        RECT 9.515 0.255 9.845 0.735 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.580 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.090 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.090 0.635 0.840 0.805 ;
        RECT 0.090 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 2.465 ;
        RECT 1.850 2.175 2.100 2.635 ;
        RECT 2.270 2.135 2.520 2.465 ;
        RECT 2.735 2.135 3.415 2.465 ;
        RECT 2.270 2.005 2.440 2.135 ;
        RECT 2.045 1.835 2.440 2.005 ;
        RECT 2.045 0.475 2.215 1.835 ;
        RECT 2.610 1.575 3.075 1.965 ;
        RECT 2.385 0.765 2.735 1.385 ;
        RECT 2.905 0.985 3.075 1.575 ;
        RECT 3.245 1.355 3.415 2.135 ;
        RECT 3.585 2.035 3.755 2.375 ;
        RECT 3.990 2.205 4.320 2.635 ;
        RECT 4.490 2.035 4.660 2.375 ;
        RECT 4.955 2.175 5.325 2.635 ;
        RECT 3.585 1.865 4.660 2.035 ;
        RECT 5.495 2.005 5.665 2.465 ;
        RECT 5.900 2.125 6.770 2.465 ;
        RECT 6.940 2.175 7.190 2.635 ;
        RECT 5.105 1.835 5.665 2.005 ;
        RECT 5.105 1.695 5.275 1.835 ;
        RECT 3.775 1.525 5.275 1.695 ;
        RECT 5.970 1.665 6.430 1.955 ;
        RECT 3.245 1.185 4.935 1.355 ;
        RECT 2.905 0.765 3.260 0.985 ;
        RECT 3.430 0.475 3.600 1.185 ;
        RECT 3.805 0.765 4.595 1.015 ;
        RECT 4.765 1.005 4.935 1.185 ;
        RECT 5.105 0.835 5.275 1.525 ;
        RECT 1.545 0.085 1.875 0.445 ;
        RECT 2.045 0.305 2.540 0.475 ;
        RECT 2.745 0.305 3.600 0.475 ;
        RECT 4.475 0.085 4.805 0.545 ;
        RECT 5.015 0.445 5.275 0.835 ;
        RECT 5.465 1.655 6.430 1.665 ;
        RECT 6.600 1.745 6.770 2.125 ;
        RECT 7.360 2.085 7.530 2.375 ;
        RECT 7.710 2.255 8.040 2.635 ;
        RECT 7.360 1.915 8.160 2.085 ;
        RECT 5.465 1.495 6.140 1.655 ;
        RECT 6.600 1.575 7.820 1.745 ;
        RECT 5.465 0.705 5.675 1.495 ;
        RECT 6.600 1.485 6.770 1.575 ;
        RECT 5.845 0.705 6.195 1.325 ;
        RECT 6.365 1.315 6.770 1.485 ;
        RECT 6.365 0.535 6.535 1.315 ;
        RECT 6.705 0.865 6.925 1.145 ;
        RECT 7.105 1.035 7.645 1.405 ;
        RECT 7.990 1.295 8.160 1.915 ;
        RECT 8.335 1.575 8.505 2.635 ;
        RECT 9.175 1.795 9.345 2.635 ;
        RECT 10.015 1.795 10.185 2.635 ;
        RECT 6.705 0.695 7.235 0.865 ;
        RECT 5.015 0.275 5.365 0.445 ;
        RECT 5.585 0.255 6.535 0.535 ;
        RECT 6.705 0.085 6.895 0.525 ;
        RECT 7.065 0.465 7.235 0.695 ;
        RECT 7.405 0.635 7.645 1.035 ;
        RECT 7.815 1.285 8.160 1.295 ;
        RECT 7.815 1.075 9.845 1.285 ;
        RECT 7.815 0.820 8.140 1.075 ;
        RECT 7.815 0.465 8.135 0.820 ;
        RECT 7.065 0.295 8.135 0.465 ;
        RECT 8.335 0.085 8.505 0.895 ;
        RECT 9.175 0.085 9.345 0.555 ;
        RECT 10.015 0.085 10.185 0.555 ;
        RECT 0.000 -0.085 10.580 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 0.610 1.105 0.780 1.275 ;
        RECT 1.015 1.785 1.185 1.955 ;
        RECT 2.905 1.785 3.075 1.955 ;
        RECT 2.445 1.105 2.615 1.275 ;
        RECT 6.025 1.785 6.195 1.955 ;
        RECT 4.165 0.765 4.335 0.935 ;
        RECT 6.025 1.105 6.195 1.275 ;
        RECT 7.105 1.080 7.275 1.250 ;
        RECT 7.405 0.765 7.575 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
      LAYER met1 ;
        RECT 0.955 1.940 1.245 1.985 ;
        RECT 2.845 1.940 3.135 1.985 ;
        RECT 5.965 1.940 6.255 1.985 ;
        RECT 0.955 1.800 6.255 1.940 ;
        RECT 0.955 1.755 1.245 1.800 ;
        RECT 2.845 1.755 3.135 1.800 ;
        RECT 5.965 1.755 6.255 1.800 ;
        RECT 0.550 1.260 0.840 1.305 ;
        RECT 2.385 1.260 2.675 1.305 ;
        RECT 5.965 1.260 6.255 1.305 ;
        RECT 0.550 1.120 6.255 1.260 ;
        RECT 0.550 1.075 0.840 1.120 ;
        RECT 2.385 1.075 2.675 1.120 ;
        RECT 5.965 1.075 6.255 1.120 ;
  END
END sky130_fd_sc_hd__dfrtp_4

#--------EOF---------

MACRO sky130_fd_sc_hd__dfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfsbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.580 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.770 1.005 2.180 1.625 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 3.765 0.920 4.055 0.965 ;
        RECT 6.985 0.920 7.275 0.965 ;
        RECT 3.765 0.780 7.275 0.920 ;
        RECT 3.765 0.735 4.055 0.780 ;
        RECT 6.985 0.735 7.275 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.580 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.365 0.785 2.285 1.005 ;
        RECT 7.860 0.905 10.205 1.015 ;
        RECT 6.930 0.785 10.205 0.905 ;
        RECT 0.005 0.105 10.205 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.770 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.580 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 9.865 1.445 10.125 2.465 ;
        RECT 9.910 0.825 10.125 1.445 ;
        RECT 9.865 0.255 10.125 0.825 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 8.370 0.255 8.700 2.465 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.580 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.175 0.635 0.840 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.240 2.465 ;
        RECT 1.455 2.135 1.785 2.635 ;
        RECT 1.955 1.965 2.125 2.465 ;
        RECT 2.360 2.250 3.190 2.420 ;
        RECT 3.430 2.255 3.810 2.635 ;
        RECT 1.430 1.795 2.125 1.965 ;
        RECT 1.430 0.825 1.600 1.795 ;
        RECT 2.350 1.575 2.850 1.955 ;
        RECT 1.430 0.635 2.125 0.825 ;
        RECT 2.350 0.705 2.570 1.575 ;
        RECT 3.020 1.405 3.190 2.250 ;
        RECT 3.990 2.085 4.160 2.375 ;
        RECT 4.330 2.255 4.660 2.635 ;
        RECT 5.110 2.165 5.760 2.415 ;
        RECT 5.930 2.255 6.340 2.635 ;
        RECT 5.590 2.085 5.760 2.165 ;
        RECT 6.540 2.085 6.780 2.375 ;
        RECT 3.360 1.835 4.710 2.085 ;
        RECT 3.360 1.575 3.610 1.835 ;
        RECT 4.120 1.405 4.370 1.565 ;
        RECT 3.020 1.235 4.370 1.405 ;
        RECT 3.020 1.195 3.440 1.235 ;
        RECT 2.750 0.645 3.100 1.015 ;
        RECT 1.455 0.085 1.785 0.465 ;
        RECT 1.955 0.305 2.125 0.635 ;
        RECT 3.270 0.465 3.440 1.195 ;
        RECT 4.540 1.065 4.710 1.835 ;
        RECT 3.610 0.735 4.020 1.065 ;
        RECT 4.310 0.725 4.710 1.065 ;
        RECT 4.900 1.655 5.400 1.965 ;
        RECT 5.590 1.915 6.780 2.085 ;
        RECT 7.010 1.945 7.340 2.635 ;
        RECT 4.900 0.895 5.070 1.655 ;
        RECT 5.240 1.065 5.420 1.475 ;
        RECT 5.590 1.405 5.760 1.915 ;
        RECT 7.510 1.765 7.680 2.375 ;
        RECT 7.510 1.745 7.830 1.765 ;
        RECT 5.930 1.575 7.830 1.745 ;
        RECT 5.590 1.235 7.470 1.405 ;
        RECT 5.820 0.895 6.150 1.015 ;
        RECT 4.900 0.725 6.150 0.895 ;
        RECT 2.425 0.265 3.440 0.465 ;
        RECT 3.610 0.085 4.020 0.525 ;
        RECT 4.310 0.295 4.560 0.725 ;
        RECT 4.740 0.085 5.080 0.545 ;
        RECT 6.320 0.475 6.490 1.235 ;
        RECT 7.140 1.175 7.470 1.235 ;
        RECT 6.660 1.005 6.990 1.065 ;
        RECT 6.660 0.735 7.320 1.005 ;
        RECT 7.640 0.680 7.830 1.575 ;
        RECT 8.020 1.480 8.200 2.635 ;
        RECT 8.890 1.325 9.220 2.465 ;
        RECT 9.445 1.825 9.615 2.635 ;
        RECT 8.890 0.995 9.740 1.325 ;
        RECT 5.640 0.305 6.490 0.475 ;
        RECT 6.670 0.085 7.330 0.565 ;
        RECT 7.510 0.350 7.830 0.680 ;
        RECT 8.020 0.085 8.200 0.905 ;
        RECT 8.890 0.255 9.220 0.995 ;
        RECT 9.445 0.085 9.615 0.585 ;
        RECT 0.000 -0.085 10.580 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 0.645 1.785 0.815 1.955 ;
        RECT 1.065 0.765 1.235 0.935 ;
        RECT 2.445 1.785 2.615 1.955 ;
        RECT 2.905 0.765 3.075 0.935 ;
        RECT 3.825 0.765 3.995 0.935 ;
        RECT 5.205 1.785 5.375 1.955 ;
        RECT 5.245 1.105 5.415 1.275 ;
        RECT 7.045 0.765 7.215 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
      LAYER met1 ;
        RECT 0.585 1.940 0.875 1.985 ;
        RECT 2.385 1.940 2.675 1.985 ;
        RECT 5.145 1.940 5.435 1.985 ;
        RECT 0.585 1.800 5.435 1.940 ;
        RECT 0.585 1.755 0.875 1.800 ;
        RECT 2.385 1.755 2.675 1.800 ;
        RECT 5.145 1.755 5.435 1.800 ;
        RECT 5.185 1.260 5.475 1.305 ;
        RECT 2.920 1.120 5.475 1.260 ;
        RECT 2.920 0.965 3.135 1.120 ;
        RECT 5.185 1.075 5.475 1.120 ;
        RECT 1.005 0.920 1.295 0.965 ;
        RECT 2.845 0.920 3.135 0.965 ;
        RECT 1.005 0.780 3.135 0.920 ;
        RECT 1.005 0.735 1.295 0.780 ;
        RECT 2.845 0.735 3.135 0.780 ;
  END
END sky130_fd_sc_hd__dfsbp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dfsbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfsbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.770 1.005 2.180 1.625 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 3.765 0.920 4.055 0.965 ;
        RECT 6.985 0.920 7.275 0.965 ;
        RECT 3.765 0.780 7.275 0.920 ;
        RECT 3.765 0.735 4.055 0.780 ;
        RECT 6.985 0.735 7.275 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.365 0.785 2.285 1.005 ;
        RECT 7.860 0.905 10.990 1.015 ;
        RECT 6.930 0.785 10.990 0.905 ;
        RECT 0.005 0.105 10.990 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 10.150 1.665 10.480 2.465 ;
        RECT 10.150 1.495 10.915 1.665 ;
        RECT 10.360 0.845 10.915 1.495 ;
        RECT 10.345 0.825 10.915 0.845 ;
        RECT 10.230 0.720 10.915 0.825 ;
        RECT 10.230 0.255 10.480 0.720 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 8.370 0.255 8.700 2.465 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.175 0.635 0.840 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.240 2.465 ;
        RECT 1.455 2.135 1.785 2.635 ;
        RECT 1.955 1.965 2.125 2.465 ;
        RECT 2.360 2.250 3.190 2.420 ;
        RECT 3.430 2.255 3.810 2.635 ;
        RECT 1.430 1.795 2.125 1.965 ;
        RECT 1.430 0.825 1.600 1.795 ;
        RECT 2.350 1.575 2.850 1.955 ;
        RECT 1.430 0.635 2.125 0.825 ;
        RECT 2.350 0.705 2.570 1.575 ;
        RECT 3.020 1.405 3.190 2.250 ;
        RECT 3.990 2.085 4.160 2.375 ;
        RECT 4.330 2.255 4.660 2.635 ;
        RECT 5.110 2.165 5.760 2.415 ;
        RECT 5.930 2.255 6.340 2.635 ;
        RECT 5.590 2.085 5.760 2.165 ;
        RECT 6.540 2.085 6.780 2.375 ;
        RECT 3.360 1.835 4.710 2.085 ;
        RECT 3.360 1.575 3.610 1.835 ;
        RECT 4.120 1.405 4.370 1.565 ;
        RECT 3.020 1.235 4.370 1.405 ;
        RECT 3.020 1.195 3.440 1.235 ;
        RECT 2.750 0.645 3.100 1.015 ;
        RECT 1.455 0.085 1.785 0.465 ;
        RECT 1.955 0.305 2.125 0.635 ;
        RECT 3.270 0.465 3.440 1.195 ;
        RECT 4.540 1.065 4.710 1.835 ;
        RECT 3.610 0.735 4.020 1.065 ;
        RECT 4.310 0.725 4.710 1.065 ;
        RECT 4.900 1.655 5.400 1.965 ;
        RECT 5.590 1.915 6.780 2.085 ;
        RECT 7.010 1.945 7.340 2.635 ;
        RECT 4.900 0.895 5.070 1.655 ;
        RECT 5.240 1.065 5.420 1.475 ;
        RECT 5.590 1.405 5.760 1.915 ;
        RECT 7.510 1.765 7.680 2.375 ;
        RECT 7.510 1.745 7.830 1.765 ;
        RECT 5.930 1.575 7.830 1.745 ;
        RECT 5.590 1.235 7.470 1.405 ;
        RECT 5.820 0.895 6.150 1.015 ;
        RECT 4.900 0.725 6.150 0.895 ;
        RECT 2.425 0.265 3.440 0.465 ;
        RECT 3.610 0.085 4.020 0.525 ;
        RECT 4.310 0.295 4.560 0.725 ;
        RECT 4.740 0.085 5.080 0.545 ;
        RECT 6.320 0.475 6.490 1.235 ;
        RECT 7.140 1.175 7.470 1.235 ;
        RECT 6.660 1.005 6.990 1.065 ;
        RECT 6.660 0.735 7.320 1.005 ;
        RECT 7.640 0.680 7.830 1.575 ;
        RECT 8.020 1.480 8.200 2.635 ;
        RECT 8.870 1.480 9.120 2.635 ;
        RECT 9.310 1.325 9.640 2.465 ;
        RECT 9.810 1.495 9.980 2.635 ;
        RECT 10.650 1.835 10.915 2.635 ;
        RECT 9.310 0.995 10.190 1.325 ;
        RECT 5.640 0.305 6.490 0.475 ;
        RECT 6.670 0.085 7.330 0.565 ;
        RECT 7.510 0.350 7.830 0.680 ;
        RECT 8.020 0.085 8.200 0.905 ;
        RECT 8.870 0.085 9.120 0.905 ;
        RECT 9.310 0.255 9.560 0.995 ;
        RECT 9.730 0.085 10.060 0.825 ;
        RECT 10.650 0.085 10.915 0.550 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 0.645 1.785 0.815 1.955 ;
        RECT 1.065 0.765 1.235 0.935 ;
        RECT 2.445 1.785 2.615 1.955 ;
        RECT 2.905 0.765 3.075 0.935 ;
        RECT 3.825 0.765 3.995 0.935 ;
        RECT 5.205 1.785 5.375 1.955 ;
        RECT 5.245 1.105 5.415 1.275 ;
        RECT 7.045 0.765 7.215 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
      LAYER met1 ;
        RECT 0.585 1.940 0.875 1.985 ;
        RECT 2.385 1.940 2.675 1.985 ;
        RECT 5.145 1.940 5.435 1.985 ;
        RECT 0.585 1.800 5.435 1.940 ;
        RECT 0.585 1.755 0.875 1.800 ;
        RECT 2.385 1.755 2.675 1.800 ;
        RECT 5.145 1.755 5.435 1.800 ;
        RECT 5.185 1.260 5.475 1.305 ;
        RECT 2.920 1.120 5.475 1.260 ;
        RECT 2.920 0.965 3.135 1.120 ;
        RECT 5.185 1.075 5.475 1.120 ;
        RECT 1.005 0.920 1.295 0.965 ;
        RECT 2.845 0.920 3.135 0.965 ;
        RECT 1.005 0.780 3.135 0.920 ;
        RECT 1.005 0.735 1.295 0.780 ;
        RECT 2.845 0.735 3.135 0.780 ;
  END
END sky130_fd_sc_hd__dfsbp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfstp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.770 1.005 2.180 1.625 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 3.790 0.920 4.080 0.965 ;
        RECT 7.050 0.920 7.340 0.965 ;
        RECT 3.790 0.780 7.340 0.920 ;
        RECT 3.790 0.735 4.080 0.780 ;
        RECT 7.050 0.735 7.340 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.365 0.785 2.285 1.005 ;
        RECT 8.365 0.905 9.285 1.015 ;
        RECT 6.950 0.785 9.285 0.905 ;
        RECT 0.005 0.105 9.285 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 8.945 1.655 9.200 2.325 ;
        RECT 9.020 0.795 9.200 1.655 ;
        RECT 8.945 0.265 9.200 0.795 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.175 0.635 0.840 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.240 2.465 ;
        RECT 1.455 2.135 1.785 2.635 ;
        RECT 1.955 1.965 2.125 2.465 ;
        RECT 2.360 2.250 3.190 2.420 ;
        RECT 3.430 2.255 3.810 2.635 ;
        RECT 1.430 1.795 2.125 1.965 ;
        RECT 1.430 0.825 1.600 1.795 ;
        RECT 2.350 1.575 2.850 1.955 ;
        RECT 1.430 0.635 2.125 0.825 ;
        RECT 2.350 0.705 2.570 1.575 ;
        RECT 3.020 1.405 3.190 2.250 ;
        RECT 3.990 2.085 4.160 2.375 ;
        RECT 4.330 2.255 4.660 2.635 ;
        RECT 5.130 2.165 5.760 2.415 ;
        RECT 5.940 2.255 6.360 2.635 ;
        RECT 5.590 2.085 5.760 2.165 ;
        RECT 6.560 2.085 6.800 2.375 ;
        RECT 3.360 1.835 4.730 2.085 ;
        RECT 3.360 1.575 3.610 1.835 ;
        RECT 4.120 1.405 4.370 1.565 ;
        RECT 3.020 1.235 4.370 1.405 ;
        RECT 3.020 1.195 3.440 1.235 ;
        RECT 2.750 0.645 3.100 1.015 ;
        RECT 1.455 0.085 1.785 0.465 ;
        RECT 1.955 0.305 2.125 0.635 ;
        RECT 3.270 0.465 3.440 1.195 ;
        RECT 4.540 1.065 4.730 1.835 ;
        RECT 3.610 0.735 4.020 1.065 ;
        RECT 4.310 0.725 4.730 1.065 ;
        RECT 4.900 1.655 5.420 1.965 ;
        RECT 5.590 1.915 6.800 2.085 ;
        RECT 7.030 1.945 7.360 2.635 ;
        RECT 4.900 0.895 5.070 1.655 ;
        RECT 5.240 1.065 5.420 1.475 ;
        RECT 5.590 1.405 5.760 1.915 ;
        RECT 7.530 1.765 7.700 2.375 ;
        RECT 7.970 1.915 8.300 2.425 ;
        RECT 7.530 1.745 7.850 1.765 ;
        RECT 5.930 1.575 7.850 1.745 ;
        RECT 5.590 1.235 7.490 1.405 ;
        RECT 5.820 0.895 6.150 1.015 ;
        RECT 4.900 0.725 6.150 0.895 ;
        RECT 2.425 0.265 3.440 0.465 ;
        RECT 3.610 0.085 4.020 0.525 ;
        RECT 4.310 0.295 4.560 0.725 ;
        RECT 4.760 0.085 5.080 0.545 ;
        RECT 6.320 0.475 6.490 1.235 ;
        RECT 7.160 1.175 7.490 1.235 ;
        RECT 6.680 1.005 7.010 1.065 ;
        RECT 6.680 0.735 7.340 1.005 ;
        RECT 7.660 0.680 7.850 1.575 ;
        RECT 5.640 0.305 6.490 0.475 ;
        RECT 6.690 0.085 7.350 0.565 ;
        RECT 7.530 0.350 7.850 0.680 ;
        RECT 8.050 1.325 8.300 1.915 ;
        RECT 8.480 1.835 8.765 2.635 ;
        RECT 8.050 0.995 8.850 1.325 ;
        RECT 8.050 0.345 8.300 0.995 ;
        RECT 8.480 0.085 8.765 0.545 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.610 1.785 0.780 1.955 ;
        RECT 1.070 0.765 1.240 0.935 ;
        RECT 2.470 1.785 2.640 1.955 ;
        RECT 2.930 0.765 3.100 0.935 ;
        RECT 3.850 0.765 4.020 0.935 ;
        RECT 5.250 1.785 5.420 1.955 ;
        RECT 5.250 1.105 5.420 1.275 ;
        RECT 7.110 0.765 7.280 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 0.550 1.940 0.840 1.985 ;
        RECT 2.410 1.940 2.700 1.985 ;
        RECT 5.190 1.940 5.480 1.985 ;
        RECT 0.550 1.800 5.480 1.940 ;
        RECT 0.550 1.755 0.840 1.800 ;
        RECT 2.410 1.755 2.700 1.800 ;
        RECT 5.190 1.755 5.480 1.800 ;
        RECT 5.190 1.260 5.480 1.305 ;
        RECT 2.945 1.120 5.480 1.260 ;
        RECT 2.945 0.965 3.160 1.120 ;
        RECT 5.190 1.075 5.480 1.120 ;
        RECT 1.010 0.920 1.300 0.965 ;
        RECT 2.870 0.920 3.160 0.965 ;
        RECT 1.010 0.780 3.160 0.920 ;
        RECT 1.010 0.735 1.300 0.780 ;
        RECT 2.870 0.735 3.160 0.780 ;
  END
END sky130_fd_sc_hd__dfstp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfstp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.770 1.005 2.180 1.625 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 3.765 0.920 4.055 0.965 ;
        RECT 6.985 0.920 7.275 0.965 ;
        RECT 3.765 0.780 7.275 0.920 ;
        RECT 3.765 0.735 4.055 0.780 ;
        RECT 6.985 0.735 7.275 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.365 0.785 2.285 1.005 ;
        RECT 7.880 0.905 9.650 1.015 ;
        RECT 6.950 0.785 9.650 0.905 ;
        RECT 0.005 0.105 9.650 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 8.810 1.615 9.140 2.460 ;
        RECT 8.810 1.495 9.575 1.615 ;
        RECT 8.975 1.445 9.575 1.495 ;
        RECT 9.020 0.895 9.575 1.445 ;
        RECT 8.990 0.855 9.575 0.895 ;
        RECT 8.975 0.825 9.575 0.855 ;
        RECT 8.890 0.765 9.575 0.825 ;
        RECT 8.890 0.265 9.135 0.765 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.085 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.015 2.045 1.235 2.465 ;
        RECT 1.455 2.135 1.785 2.635 ;
        RECT 0.085 1.795 0.835 1.965 ;
        RECT 0.605 0.805 0.835 1.795 ;
        RECT 0.085 0.635 0.835 0.805 ;
        RECT 0.085 0.345 0.345 0.635 ;
        RECT 1.005 0.565 1.235 2.045 ;
        RECT 1.955 1.965 2.125 2.465 ;
        RECT 2.360 2.250 3.190 2.420 ;
        RECT 3.430 2.255 3.810 2.635 ;
        RECT 1.430 1.795 2.125 1.965 ;
        RECT 1.430 0.825 1.600 1.795 ;
        RECT 2.350 1.575 2.850 1.955 ;
        RECT 1.430 0.635 2.125 0.825 ;
        RECT 2.350 0.705 2.570 1.575 ;
        RECT 3.020 1.405 3.190 2.250 ;
        RECT 3.990 2.085 4.160 2.375 ;
        RECT 4.330 2.255 4.660 2.635 ;
        RECT 5.110 2.165 5.740 2.415 ;
        RECT 5.920 2.255 6.340 2.635 ;
        RECT 5.570 2.085 5.740 2.165 ;
        RECT 6.540 2.085 6.780 2.375 ;
        RECT 3.360 1.835 4.710 2.085 ;
        RECT 3.360 1.575 3.610 1.835 ;
        RECT 4.120 1.405 4.370 1.565 ;
        RECT 3.020 1.235 4.370 1.405 ;
        RECT 3.020 1.195 3.440 1.235 ;
        RECT 2.750 0.645 3.100 1.015 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.235 0.565 ;
        RECT 1.455 0.085 1.785 0.465 ;
        RECT 1.955 0.305 2.125 0.635 ;
        RECT 3.270 0.465 3.440 1.195 ;
        RECT 4.540 1.065 4.710 1.835 ;
        RECT 3.610 0.735 4.020 1.065 ;
        RECT 4.310 0.725 4.710 1.065 ;
        RECT 4.880 1.655 5.400 1.965 ;
        RECT 5.570 1.915 6.780 2.085 ;
        RECT 7.010 1.945 7.340 2.635 ;
        RECT 4.880 0.895 5.050 1.655 ;
        RECT 5.220 1.065 5.400 1.475 ;
        RECT 5.570 1.405 5.740 1.915 ;
        RECT 7.510 1.765 7.680 2.375 ;
        RECT 7.970 1.915 8.300 2.425 ;
        RECT 7.510 1.745 7.880 1.765 ;
        RECT 5.910 1.575 7.880 1.745 ;
        RECT 5.570 1.235 7.490 1.405 ;
        RECT 5.800 0.895 6.150 1.015 ;
        RECT 4.880 0.725 6.150 0.895 ;
        RECT 2.425 0.265 3.440 0.465 ;
        RECT 3.610 0.085 4.020 0.525 ;
        RECT 4.310 0.295 4.560 0.725 ;
        RECT 4.760 0.085 5.080 0.545 ;
        RECT 6.320 0.475 6.490 1.235 ;
        RECT 7.140 1.175 7.490 1.235 ;
        RECT 6.660 1.005 7.010 1.065 ;
        RECT 6.660 0.735 7.340 1.005 ;
        RECT 7.690 0.680 7.880 1.575 ;
        RECT 5.640 0.305 6.490 0.475 ;
        RECT 6.690 0.085 7.330 0.565 ;
        RECT 7.530 0.350 7.880 0.680 ;
        RECT 8.050 1.325 8.300 1.915 ;
        RECT 8.470 1.495 8.640 2.635 ;
        RECT 9.310 1.785 9.575 2.635 ;
        RECT 8.050 0.995 8.850 1.325 ;
        RECT 8.050 0.345 8.220 0.995 ;
        RECT 8.390 0.085 8.720 0.825 ;
        RECT 9.305 0.085 9.575 0.595 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.605 1.785 0.775 1.955 ;
        RECT 1.065 0.765 1.235 0.935 ;
        RECT 2.445 1.785 2.615 1.955 ;
        RECT 2.905 0.765 3.075 0.935 ;
        RECT 3.825 0.765 3.995 0.935 ;
        RECT 5.205 1.785 5.375 1.955 ;
        RECT 5.225 1.105 5.395 1.275 ;
        RECT 7.045 0.765 7.215 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 0.545 1.940 0.835 1.985 ;
        RECT 2.385 1.940 2.675 1.985 ;
        RECT 5.145 1.940 5.435 1.985 ;
        RECT 0.545 1.800 5.435 1.940 ;
        RECT 0.545 1.755 0.835 1.800 ;
        RECT 2.385 1.755 2.675 1.800 ;
        RECT 5.145 1.755 5.435 1.800 ;
        RECT 5.165 1.260 5.455 1.305 ;
        RECT 2.920 1.120 5.455 1.260 ;
        RECT 2.920 0.965 3.135 1.120 ;
        RECT 5.165 1.075 5.455 1.120 ;
        RECT 1.005 0.920 1.295 0.965 ;
        RECT 2.845 0.920 3.135 0.965 ;
        RECT 1.005 0.780 3.135 0.920 ;
        RECT 1.005 0.735 1.295 0.780 ;
        RECT 2.845 0.735 3.135 0.780 ;
  END
END sky130_fd_sc_hd__dfstp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dfstp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfstp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 1.770 1.005 2.180 1.625 ;
    END
  END D
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 3.765 0.920 4.055 0.965 ;
        RECT 6.985 0.920 7.275 0.965 ;
        RECT 3.765 0.780 7.275 0.920 ;
        RECT 3.765 0.735 4.055 0.780 ;
        RECT 6.985 0.735 7.275 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.365 0.785 2.285 1.005 ;
        RECT 8.345 0.905 10.945 1.015 ;
        RECT 6.930 0.785 10.945 0.905 ;
        RECT 0.005 0.105 10.945 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.320000 ;
    PORT
      LAYER li1 ;
        RECT 8.925 1.640 9.170 2.465 ;
        RECT 9.765 1.640 9.935 2.465 ;
        RECT 10.605 1.640 10.955 2.465 ;
        RECT 8.925 1.470 10.955 1.640 ;
        RECT 10.725 0.885 10.955 1.470 ;
        RECT 8.925 0.715 10.955 0.885 ;
        RECT 8.925 0.265 9.170 0.715 ;
        RECT 9.765 0.265 9.935 0.715 ;
        RECT 10.605 0.265 10.955 0.715 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.175 0.635 0.840 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.240 2.465 ;
        RECT 1.455 2.135 1.785 2.635 ;
        RECT 1.955 1.965 2.125 2.465 ;
        RECT 2.360 2.250 3.190 2.420 ;
        RECT 3.430 2.255 3.810 2.635 ;
        RECT 1.430 1.795 2.125 1.965 ;
        RECT 1.430 0.825 1.600 1.795 ;
        RECT 2.350 1.575 2.850 1.955 ;
        RECT 1.430 0.635 2.125 0.825 ;
        RECT 2.350 0.705 2.570 1.575 ;
        RECT 3.020 1.405 3.190 2.250 ;
        RECT 3.990 2.085 4.160 2.375 ;
        RECT 4.330 2.255 4.660 2.635 ;
        RECT 5.110 2.165 5.740 2.415 ;
        RECT 5.920 2.255 6.340 2.635 ;
        RECT 5.570 2.085 5.740 2.165 ;
        RECT 6.540 2.085 6.780 2.375 ;
        RECT 3.360 1.835 4.710 2.085 ;
        RECT 3.360 1.575 3.610 1.835 ;
        RECT 4.120 1.405 4.370 1.565 ;
        RECT 3.020 1.235 4.370 1.405 ;
        RECT 3.020 1.195 3.440 1.235 ;
        RECT 2.750 0.645 3.100 1.015 ;
        RECT 1.455 0.085 1.785 0.465 ;
        RECT 1.955 0.305 2.125 0.635 ;
        RECT 3.270 0.465 3.440 1.195 ;
        RECT 4.540 1.065 4.710 1.835 ;
        RECT 3.610 0.735 4.020 1.065 ;
        RECT 4.310 0.725 4.710 1.065 ;
        RECT 4.880 1.655 5.400 1.965 ;
        RECT 5.570 1.915 6.780 2.085 ;
        RECT 7.010 1.945 7.340 2.635 ;
        RECT 4.880 0.895 5.050 1.655 ;
        RECT 5.220 1.065 5.400 1.475 ;
        RECT 5.570 1.405 5.740 1.915 ;
        RECT 7.510 1.765 7.680 2.375 ;
        RECT 7.950 1.915 8.280 2.425 ;
        RECT 7.510 1.745 7.850 1.765 ;
        RECT 5.910 1.575 7.850 1.745 ;
        RECT 5.570 1.235 7.470 1.405 ;
        RECT 5.820 0.895 6.150 1.015 ;
        RECT 4.880 0.725 6.150 0.895 ;
        RECT 2.425 0.265 3.440 0.465 ;
        RECT 3.610 0.085 4.020 0.525 ;
        RECT 4.310 0.295 4.560 0.725 ;
        RECT 4.740 0.085 5.080 0.545 ;
        RECT 6.320 0.475 6.490 1.235 ;
        RECT 7.140 1.175 7.470 1.235 ;
        RECT 6.660 1.005 6.990 1.065 ;
        RECT 6.660 0.735 7.320 1.005 ;
        RECT 7.640 0.680 7.850 1.575 ;
        RECT 5.640 0.305 6.490 0.475 ;
        RECT 6.670 0.085 7.330 0.565 ;
        RECT 7.510 0.350 7.850 0.680 ;
        RECT 8.030 1.275 8.280 1.915 ;
        RECT 8.460 1.835 8.745 2.635 ;
        RECT 9.340 1.810 9.595 2.635 ;
        RECT 10.105 1.810 10.435 2.635 ;
        RECT 8.030 1.055 10.555 1.275 ;
        RECT 8.030 0.345 8.280 1.055 ;
        RECT 8.460 0.085 8.745 0.545 ;
        RECT 9.340 0.085 9.595 0.545 ;
        RECT 10.105 0.085 10.435 0.545 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 0.615 1.785 0.785 1.955 ;
        RECT 1.065 0.765 1.235 0.935 ;
        RECT 2.445 1.785 2.615 1.955 ;
        RECT 2.905 0.765 3.075 0.935 ;
        RECT 3.825 0.765 3.995 0.935 ;
        RECT 5.205 1.785 5.375 1.955 ;
        RECT 5.225 1.105 5.395 1.275 ;
        RECT 7.045 0.765 7.215 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
      LAYER met1 ;
        RECT 0.555 1.940 0.845 1.985 ;
        RECT 2.385 1.940 2.675 1.985 ;
        RECT 5.145 1.940 5.435 1.985 ;
        RECT 0.555 1.800 5.435 1.940 ;
        RECT 0.555 1.755 0.845 1.800 ;
        RECT 2.385 1.755 2.675 1.800 ;
        RECT 5.145 1.755 5.435 1.800 ;
        RECT 5.165 1.260 5.455 1.305 ;
        RECT 2.920 1.120 5.455 1.260 ;
        RECT 2.920 0.965 3.135 1.120 ;
        RECT 5.165 1.075 5.455 1.120 ;
        RECT 1.005 0.920 1.295 0.965 ;
        RECT 2.845 0.920 3.135 0.965 ;
        RECT 1.005 0.780 3.135 0.920 ;
        RECT 1.005 0.735 1.295 0.780 ;
        RECT 2.845 0.735 3.135 0.780 ;
  END
END sky130_fd_sc_hd__dfstp_4

#--------EOF---------

MACRO sky130_fd_sc_hd__dfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.370 0.715 1.650 1.665 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.520 0.785 4.430 1.005 ;
        RECT 5.970 0.785 8.735 1.015 ;
        RECT 0.005 0.105 8.735 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 6.890 1.575 7.220 2.420 ;
        RECT 6.890 1.495 7.300 1.575 ;
        RECT 7.065 1.445 7.300 1.495 ;
        RECT 7.110 0.865 7.300 1.445 ;
        RECT 7.055 0.825 7.300 0.865 ;
        RECT 6.900 0.740 7.300 0.825 ;
        RECT 6.900 0.305 7.230 0.740 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 8.315 1.480 8.650 2.465 ;
        RECT 8.415 0.910 8.650 1.480 ;
        RECT 8.395 0.255 8.650 0.910 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.740 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.175 0.635 0.840 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.200 2.465 ;
        RECT 1.440 2.175 1.705 2.635 ;
        RECT 1.875 2.040 2.125 2.465 ;
        RECT 2.335 2.190 3.440 2.360 ;
        RECT 1.820 1.910 2.125 2.040 ;
        RECT 1.820 0.805 1.990 1.910 ;
        RECT 2.160 1.125 2.400 1.720 ;
        RECT 2.570 1.655 3.100 2.020 ;
        RECT 2.570 0.955 2.740 1.655 ;
        RECT 3.270 1.575 3.440 2.190 ;
        RECT 3.610 1.835 3.780 2.635 ;
        RECT 3.950 2.135 4.200 2.465 ;
        RECT 4.425 2.165 5.310 2.335 ;
        RECT 3.270 1.485 3.780 1.575 ;
        RECT 1.820 0.675 2.045 0.805 ;
        RECT 2.215 0.735 2.740 0.955 ;
        RECT 2.910 1.315 3.780 1.485 ;
        RECT 1.455 0.085 1.705 0.545 ;
        RECT 1.875 0.535 2.045 0.675 ;
        RECT 2.910 0.535 3.080 1.315 ;
        RECT 3.610 1.245 3.780 1.315 ;
        RECT 3.290 1.065 3.490 1.095 ;
        RECT 3.950 1.065 4.120 2.135 ;
        RECT 4.290 1.245 4.480 1.965 ;
        RECT 3.290 0.765 4.120 1.065 ;
        RECT 4.650 1.035 4.970 1.995 ;
        RECT 1.875 0.365 2.210 0.535 ;
        RECT 2.405 0.365 3.080 0.535 ;
        RECT 3.400 0.085 3.770 0.585 ;
        RECT 3.950 0.535 4.120 0.765 ;
        RECT 4.505 0.705 4.970 1.035 ;
        RECT 5.140 1.325 5.310 2.165 ;
        RECT 5.490 2.135 5.805 2.635 ;
        RECT 6.040 1.905 6.380 2.465 ;
        RECT 5.480 1.530 6.380 1.905 ;
        RECT 6.550 1.625 6.720 2.635 ;
        RECT 7.410 1.715 7.740 2.445 ;
        RECT 6.190 1.325 6.380 1.530 ;
        RECT 7.470 1.325 7.740 1.715 ;
        RECT 7.930 1.495 8.145 2.635 ;
        RECT 5.140 0.995 6.020 1.325 ;
        RECT 6.190 0.995 6.940 1.325 ;
        RECT 7.470 0.995 8.245 1.325 ;
        RECT 5.140 0.535 5.310 0.995 ;
        RECT 6.190 0.825 6.390 0.995 ;
        RECT 3.950 0.365 4.355 0.535 ;
        RECT 4.525 0.365 5.310 0.535 ;
        RECT 5.585 0.085 5.795 0.615 ;
        RECT 6.060 0.300 6.390 0.825 ;
        RECT 6.560 0.085 6.730 0.695 ;
        RECT 7.470 0.615 7.670 0.995 ;
        RECT 7.420 0.345 7.670 0.615 ;
        RECT 7.905 0.085 8.225 0.545 ;
        RECT 0.000 -0.085 8.740 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 0.630 1.785 0.800 1.955 ;
        RECT 1.025 1.445 1.195 1.615 ;
        RECT 2.730 1.785 2.900 1.955 ;
        RECT 2.215 1.445 2.385 1.615 ;
        RECT 4.300 1.785 4.470 1.955 ;
        RECT 4.735 1.445 4.905 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
      LAYER met1 ;
        RECT 0.570 1.940 0.860 1.985 ;
        RECT 2.670 1.940 2.960 1.985 ;
        RECT 4.240 1.940 4.530 1.985 ;
        RECT 0.570 1.800 4.530 1.940 ;
        RECT 0.570 1.755 0.860 1.800 ;
        RECT 2.670 1.755 2.960 1.800 ;
        RECT 4.240 1.755 4.530 1.800 ;
        RECT 0.965 1.600 1.255 1.645 ;
        RECT 2.155 1.600 2.445 1.645 ;
        RECT 4.675 1.600 4.965 1.645 ;
        RECT 0.965 1.460 4.965 1.600 ;
        RECT 0.965 1.415 1.255 1.460 ;
        RECT 2.155 1.415 2.445 1.460 ;
        RECT 4.675 1.415 4.965 1.460 ;
  END
END sky130_fd_sc_hd__dfxbp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.370 0.715 1.650 1.665 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.520 0.785 4.430 1.005 ;
        RECT 5.970 0.785 9.655 1.015 ;
        RECT 0.005 0.105 9.655 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 6.890 1.575 7.220 2.420 ;
        RECT 6.890 1.495 7.300 1.575 ;
        RECT 7.065 1.445 7.300 1.495 ;
        RECT 7.110 0.865 7.300 1.445 ;
        RECT 7.055 0.825 7.300 0.865 ;
        RECT 6.900 0.740 7.300 0.825 ;
        RECT 6.900 0.305 7.230 0.740 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 8.810 1.495 9.145 2.465 ;
        RECT 8.930 0.885 9.145 1.495 ;
        RECT 8.890 0.265 9.145 0.885 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.175 0.635 0.840 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.200 2.465 ;
        RECT 1.440 2.175 1.705 2.635 ;
        RECT 1.875 2.040 2.125 2.465 ;
        RECT 2.335 2.190 3.440 2.360 ;
        RECT 1.820 1.910 2.125 2.040 ;
        RECT 1.820 0.805 1.990 1.910 ;
        RECT 2.160 1.125 2.400 1.720 ;
        RECT 2.570 1.655 3.100 2.020 ;
        RECT 2.570 0.955 2.740 1.655 ;
        RECT 3.270 1.575 3.440 2.190 ;
        RECT 3.610 1.835 3.780 2.635 ;
        RECT 3.950 2.135 4.200 2.465 ;
        RECT 4.425 2.165 5.310 2.335 ;
        RECT 3.270 1.485 3.780 1.575 ;
        RECT 1.820 0.675 2.045 0.805 ;
        RECT 2.215 0.735 2.740 0.955 ;
        RECT 2.910 1.315 3.780 1.485 ;
        RECT 1.455 0.085 1.705 0.545 ;
        RECT 1.875 0.535 2.045 0.675 ;
        RECT 2.910 0.535 3.080 1.315 ;
        RECT 3.610 1.245 3.780 1.315 ;
        RECT 3.290 1.065 3.490 1.095 ;
        RECT 3.950 1.065 4.120 2.135 ;
        RECT 4.290 1.245 4.480 1.965 ;
        RECT 3.290 0.765 4.120 1.065 ;
        RECT 4.650 1.035 4.970 1.995 ;
        RECT 1.875 0.365 2.210 0.535 ;
        RECT 2.405 0.365 3.080 0.535 ;
        RECT 3.400 0.085 3.770 0.585 ;
        RECT 3.950 0.535 4.120 0.765 ;
        RECT 4.505 0.705 4.970 1.035 ;
        RECT 5.140 1.325 5.310 2.165 ;
        RECT 5.490 2.135 5.805 2.635 ;
        RECT 6.040 1.905 6.380 2.465 ;
        RECT 5.480 1.530 6.380 1.905 ;
        RECT 6.550 1.625 6.720 2.635 ;
        RECT 7.390 1.720 7.565 2.635 ;
        RECT 7.905 1.715 8.235 2.445 ;
        RECT 6.190 1.325 6.380 1.530 ;
        RECT 7.965 1.325 8.235 1.715 ;
        RECT 8.425 1.495 8.640 2.635 ;
        RECT 9.315 1.495 9.565 2.635 ;
        RECT 5.140 0.995 6.020 1.325 ;
        RECT 6.190 0.995 6.940 1.325 ;
        RECT 7.965 0.995 8.760 1.325 ;
        RECT 5.140 0.535 5.310 0.995 ;
        RECT 6.190 0.825 6.390 0.995 ;
        RECT 3.950 0.365 4.355 0.535 ;
        RECT 4.525 0.365 5.310 0.535 ;
        RECT 5.585 0.085 5.795 0.615 ;
        RECT 6.060 0.300 6.390 0.825 ;
        RECT 6.560 0.085 6.730 0.695 ;
        RECT 7.965 0.615 8.165 0.995 ;
        RECT 7.400 0.085 7.570 0.600 ;
        RECT 7.905 0.345 8.165 0.615 ;
        RECT 8.390 0.085 8.720 0.825 ;
        RECT 9.315 0.085 9.565 0.905 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.630 1.785 0.800 1.955 ;
        RECT 1.025 1.445 1.195 1.615 ;
        RECT 2.730 1.785 2.900 1.955 ;
        RECT 2.215 1.445 2.385 1.615 ;
        RECT 4.300 1.785 4.470 1.955 ;
        RECT 4.735 1.445 4.905 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 0.570 1.940 0.860 1.985 ;
        RECT 2.670 1.940 2.960 1.985 ;
        RECT 4.240 1.940 4.530 1.985 ;
        RECT 0.570 1.800 4.530 1.940 ;
        RECT 0.570 1.755 0.860 1.800 ;
        RECT 2.670 1.755 2.960 1.800 ;
        RECT 4.240 1.755 4.530 1.800 ;
        RECT 0.965 1.600 1.255 1.645 ;
        RECT 2.155 1.600 2.445 1.645 ;
        RECT 4.675 1.600 4.965 1.645 ;
        RECT 0.965 1.460 4.965 1.600 ;
        RECT 0.965 1.415 1.255 1.460 ;
        RECT 2.155 1.415 2.445 1.460 ;
        RECT 4.675 1.415 4.965 1.460 ;
  END
END sky130_fd_sc_hd__dfxbp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.370 0.715 1.650 1.665 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.520 0.785 4.430 1.005 ;
        RECT 5.965 0.785 7.315 1.015 ;
        RECT 0.005 0.105 7.315 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 6.885 1.575 7.215 2.420 ;
        RECT 6.885 1.495 7.275 1.575 ;
        RECT 7.060 1.445 7.275 1.495 ;
        RECT 7.105 0.865 7.275 1.445 ;
        RECT 7.050 0.825 7.275 0.865 ;
        RECT 6.895 0.740 7.275 0.825 ;
        RECT 6.895 0.305 7.225 0.740 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.175 0.635 0.840 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.200 2.465 ;
        RECT 1.440 2.175 1.705 2.635 ;
        RECT 1.875 2.040 2.125 2.465 ;
        RECT 2.335 2.190 3.440 2.360 ;
        RECT 1.820 1.910 2.125 2.040 ;
        RECT 1.820 0.805 1.990 1.910 ;
        RECT 2.160 1.125 2.400 1.720 ;
        RECT 2.570 1.655 3.100 2.020 ;
        RECT 2.570 0.955 2.740 1.655 ;
        RECT 3.270 1.575 3.440 2.190 ;
        RECT 3.610 1.835 3.780 2.635 ;
        RECT 3.950 2.135 4.200 2.465 ;
        RECT 4.425 2.165 5.310 2.335 ;
        RECT 3.270 1.485 3.780 1.575 ;
        RECT 1.820 0.675 2.045 0.805 ;
        RECT 2.215 0.735 2.740 0.955 ;
        RECT 2.910 1.315 3.780 1.485 ;
        RECT 1.455 0.085 1.705 0.545 ;
        RECT 1.875 0.535 2.045 0.675 ;
        RECT 2.910 0.535 3.080 1.315 ;
        RECT 3.610 1.245 3.780 1.315 ;
        RECT 3.290 1.065 3.490 1.095 ;
        RECT 3.950 1.065 4.120 2.135 ;
        RECT 4.290 1.245 4.480 1.965 ;
        RECT 3.290 0.765 4.120 1.065 ;
        RECT 4.650 1.035 4.970 1.995 ;
        RECT 1.875 0.365 2.210 0.535 ;
        RECT 2.405 0.365 3.080 0.535 ;
        RECT 3.400 0.085 3.770 0.585 ;
        RECT 3.950 0.535 4.120 0.765 ;
        RECT 4.505 0.705 4.970 1.035 ;
        RECT 5.140 1.325 5.310 2.165 ;
        RECT 5.490 2.135 5.805 2.635 ;
        RECT 6.035 1.905 6.375 2.465 ;
        RECT 5.480 1.530 6.375 1.905 ;
        RECT 6.545 1.625 6.715 2.635 ;
        RECT 6.185 1.325 6.375 1.530 ;
        RECT 5.140 0.995 6.015 1.325 ;
        RECT 6.185 0.995 6.935 1.325 ;
        RECT 5.140 0.535 5.310 0.995 ;
        RECT 6.185 0.825 6.385 0.995 ;
        RECT 3.950 0.365 4.355 0.535 ;
        RECT 4.525 0.365 5.310 0.535 ;
        RECT 5.585 0.085 5.795 0.615 ;
        RECT 6.055 0.300 6.385 0.825 ;
        RECT 6.555 0.085 6.725 0.695 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.630 1.785 0.800 1.955 ;
        RECT 1.025 1.445 1.195 1.615 ;
        RECT 2.730 1.785 2.900 1.955 ;
        RECT 2.215 1.445 2.385 1.615 ;
        RECT 4.300 1.785 4.470 1.955 ;
        RECT 4.735 1.445 4.905 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
      LAYER met1 ;
        RECT 0.570 1.940 0.860 1.985 ;
        RECT 2.670 1.940 2.960 1.985 ;
        RECT 4.240 1.940 4.530 1.985 ;
        RECT 0.570 1.800 4.530 1.940 ;
        RECT 0.570 1.755 0.860 1.800 ;
        RECT 2.670 1.755 2.960 1.800 ;
        RECT 4.240 1.755 4.530 1.800 ;
        RECT 0.965 1.600 1.255 1.645 ;
        RECT 2.155 1.600 2.445 1.645 ;
        RECT 4.675 1.600 4.965 1.645 ;
        RECT 0.965 1.460 4.965 1.600 ;
        RECT 0.965 1.415 1.255 1.460 ;
        RECT 2.155 1.415 2.445 1.460 ;
        RECT 4.675 1.415 4.965 1.460 ;
  END
END sky130_fd_sc_hd__dfxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.370 0.715 1.650 1.665 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.520 0.785 4.430 1.005 ;
        RECT 5.965 0.785 7.735 1.015 ;
        RECT 0.005 0.105 7.735 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 6.885 1.575 7.215 2.420 ;
        RECT 6.885 1.495 7.275 1.575 ;
        RECT 7.060 1.445 7.275 1.495 ;
        RECT 7.105 0.865 7.275 1.445 ;
        RECT 7.050 0.825 7.275 0.865 ;
        RECT 6.895 0.740 7.275 0.825 ;
        RECT 6.895 0.305 7.225 0.740 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.175 0.635 0.840 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.200 2.465 ;
        RECT 1.440 2.175 1.705 2.635 ;
        RECT 1.875 2.040 2.125 2.465 ;
        RECT 2.335 2.190 3.440 2.360 ;
        RECT 1.820 1.910 2.125 2.040 ;
        RECT 1.820 0.805 1.990 1.910 ;
        RECT 2.160 1.125 2.400 1.720 ;
        RECT 2.570 1.655 3.100 2.020 ;
        RECT 2.570 0.955 2.740 1.655 ;
        RECT 3.270 1.575 3.440 2.190 ;
        RECT 3.610 1.835 3.780 2.635 ;
        RECT 3.950 2.135 4.200 2.465 ;
        RECT 4.425 2.165 5.310 2.335 ;
        RECT 3.270 1.485 3.780 1.575 ;
        RECT 1.820 0.675 2.045 0.805 ;
        RECT 2.215 0.735 2.740 0.955 ;
        RECT 2.910 1.315 3.780 1.485 ;
        RECT 1.455 0.085 1.705 0.545 ;
        RECT 1.875 0.535 2.045 0.675 ;
        RECT 2.910 0.535 3.080 1.315 ;
        RECT 3.610 1.245 3.780 1.315 ;
        RECT 3.290 1.065 3.490 1.095 ;
        RECT 3.950 1.065 4.120 2.135 ;
        RECT 4.290 1.245 4.480 1.965 ;
        RECT 3.290 0.765 4.120 1.065 ;
        RECT 4.650 1.035 4.970 1.995 ;
        RECT 1.875 0.365 2.210 0.535 ;
        RECT 2.405 0.365 3.080 0.535 ;
        RECT 3.400 0.085 3.770 0.585 ;
        RECT 3.950 0.535 4.120 0.765 ;
        RECT 4.505 0.705 4.970 1.035 ;
        RECT 5.140 1.325 5.310 2.165 ;
        RECT 5.490 2.135 5.805 2.635 ;
        RECT 6.035 1.905 6.375 2.465 ;
        RECT 5.480 1.530 6.375 1.905 ;
        RECT 6.545 1.625 6.715 2.635 ;
        RECT 7.385 1.720 7.555 2.635 ;
        RECT 6.185 1.325 6.375 1.530 ;
        RECT 5.140 0.995 6.015 1.325 ;
        RECT 6.185 0.995 6.935 1.325 ;
        RECT 5.140 0.535 5.310 0.995 ;
        RECT 6.185 0.825 6.385 0.995 ;
        RECT 3.950 0.365 4.355 0.535 ;
        RECT 4.525 0.365 5.310 0.535 ;
        RECT 5.585 0.085 5.795 0.615 ;
        RECT 6.055 0.300 6.385 0.825 ;
        RECT 6.555 0.085 6.725 0.695 ;
        RECT 7.395 0.085 7.565 0.600 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.630 1.785 0.800 1.955 ;
        RECT 1.025 1.445 1.195 1.615 ;
        RECT 2.730 1.785 2.900 1.955 ;
        RECT 2.215 1.445 2.385 1.615 ;
        RECT 4.300 1.785 4.470 1.955 ;
        RECT 4.735 1.445 4.905 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
      LAYER met1 ;
        RECT 0.570 1.940 0.860 1.985 ;
        RECT 2.670 1.940 2.960 1.985 ;
        RECT 4.240 1.940 4.530 1.985 ;
        RECT 0.570 1.800 4.530 1.940 ;
        RECT 0.570 1.755 0.860 1.800 ;
        RECT 2.670 1.755 2.960 1.800 ;
        RECT 4.240 1.755 4.530 1.800 ;
        RECT 0.965 1.600 1.255 1.645 ;
        RECT 2.155 1.600 2.445 1.645 ;
        RECT 4.675 1.600 4.965 1.645 ;
        RECT 0.965 1.460 4.965 1.600 ;
        RECT 0.965 1.415 1.255 1.460 ;
        RECT 2.155 1.415 2.445 1.460 ;
        RECT 4.675 1.415 4.965 1.460 ;
  END
END sky130_fd_sc_hd__dfxtp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dfxtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.975 0.440 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.440 1.065 1.720 1.665 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.550 0.785 4.460 1.005 ;
        RECT 6.000 0.785 8.705 1.015 ;
        RECT 0.005 0.105 8.705 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 6.985 1.635 7.320 2.395 ;
        RECT 7.840 1.635 8.170 2.395 ;
        RECT 6.985 1.465 8.655 1.635 ;
        RECT 8.410 0.900 8.655 1.465 ;
        RECT 6.985 0.730 8.655 0.900 ;
        RECT 6.985 0.305 7.320 0.730 ;
        RECT 7.840 0.305 8.175 0.730 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.740 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.840 1.965 ;
        RECT 0.610 0.805 0.840 1.795 ;
        RECT 0.175 0.635 0.840 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.240 2.465 ;
        RECT 1.440 2.175 1.705 2.635 ;
        RECT 1.890 2.065 2.125 2.440 ;
        RECT 2.370 2.190 3.440 2.360 ;
        RECT 1.455 0.085 1.705 0.545 ;
        RECT 1.890 0.535 2.060 2.065 ;
        RECT 2.230 1.035 2.470 1.905 ;
        RECT 2.660 1.655 3.100 2.010 ;
        RECT 3.270 1.575 3.440 2.190 ;
        RECT 3.610 1.835 3.780 2.635 ;
        RECT 3.950 2.135 4.200 2.465 ;
        RECT 4.425 2.165 5.310 2.335 ;
        RECT 3.270 1.485 3.780 1.575 ;
        RECT 2.980 1.315 3.780 1.485 ;
        RECT 2.230 0.705 2.810 1.035 ;
        RECT 2.980 0.535 3.150 1.315 ;
        RECT 3.610 1.245 3.780 1.315 ;
        RECT 3.320 1.065 3.490 1.095 ;
        RECT 3.950 1.065 4.120 2.135 ;
        RECT 4.290 1.245 4.480 1.965 ;
        RECT 4.650 1.575 4.970 1.905 ;
        RECT 3.320 0.765 4.120 1.065 ;
        RECT 4.650 1.035 4.840 1.575 ;
        RECT 1.890 0.365 2.220 0.535 ;
        RECT 2.400 0.365 3.150 0.535 ;
        RECT 3.400 0.085 3.770 0.585 ;
        RECT 3.950 0.535 4.120 0.765 ;
        RECT 4.290 0.705 4.840 1.035 ;
        RECT 5.140 1.245 5.310 2.165 ;
        RECT 5.490 2.135 5.705 2.635 ;
        RECT 6.170 1.830 6.340 2.455 ;
        RECT 6.625 1.855 6.805 2.635 ;
        RECT 5.480 1.670 6.340 1.830 ;
        RECT 7.500 1.805 7.670 2.635 ;
        RECT 8.340 1.805 8.510 2.635 ;
        RECT 5.480 1.500 6.590 1.670 ;
        RECT 6.420 1.245 6.590 1.500 ;
        RECT 5.140 1.075 6.230 1.245 ;
        RECT 6.420 1.075 8.240 1.245 ;
        RECT 5.140 0.535 5.310 1.075 ;
        RECT 6.420 0.905 6.590 1.075 ;
        RECT 6.090 0.735 6.590 0.905 ;
        RECT 3.950 0.365 4.410 0.535 ;
        RECT 4.640 0.365 5.310 0.535 ;
        RECT 5.625 0.085 5.795 0.615 ;
        RECT 6.090 0.295 6.450 0.735 ;
        RECT 6.625 0.085 6.795 0.565 ;
        RECT 7.495 0.085 7.665 0.560 ;
        RECT 8.345 0.085 8.515 0.560 ;
        RECT 0.000 -0.085 8.740 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 0.610 1.785 0.780 1.955 ;
        RECT 1.070 0.765 1.240 0.935 ;
        RECT 2.930 1.785 3.100 1.955 ;
        RECT 2.470 0.765 2.640 0.935 ;
        RECT 4.310 1.785 4.480 1.955 ;
        RECT 4.310 0.765 4.480 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
      LAYER met1 ;
        RECT 0.550 1.940 0.840 1.985 ;
        RECT 2.870 1.940 3.160 1.985 ;
        RECT 4.250 1.940 4.540 1.985 ;
        RECT 0.550 1.800 4.540 1.940 ;
        RECT 0.550 1.755 0.840 1.800 ;
        RECT 2.870 1.755 3.160 1.800 ;
        RECT 4.250 1.755 4.540 1.800 ;
        RECT 1.010 0.920 1.300 0.965 ;
        RECT 2.410 0.920 2.700 0.965 ;
        RECT 4.250 0.920 4.540 0.965 ;
        RECT 1.010 0.780 4.540 0.920 ;
        RECT 1.010 0.735 1.300 0.780 ;
        RECT 2.410 0.735 2.700 0.780 ;
        RECT 4.250 0.735 4.540 0.780 ;
  END
END sky130_fd_sc_hd__dfxtp_4

#--------EOF---------

MACRO sky130_fd_sc_hd__diode_2
  CLASS CORE ANTENNACELL ;
  FOREIGN sky130_fd_sc_hd__diode_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.920 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN DIODE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.255 0.835 2.465 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 0.920 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.065 0.915 1.015 ;
        RECT 0.145 -0.085 0.315 0.065 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.110 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.920 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.920 2.805 ;
        RECT 0.000 -0.085 0.920 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
  END
END sky130_fd_sc_hd__diode_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlclkp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER met1 ;
        RECT 0.085 1.260 0.380 1.305 ;
        RECT 5.150 1.260 5.440 1.305 ;
        RECT 0.085 1.120 5.440 1.260 ;
        RECT 0.085 1.075 0.380 1.120 ;
        RECT 5.150 1.075 5.440 1.120 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.435 2.185 1.685 ;
        RECT 1.985 0.385 2.185 1.435 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.395 0.880 2.435 1.145 ;
        RECT 3.675 0.880 4.660 1.015 ;
        RECT 1.395 0.785 4.660 0.880 ;
        RECT 5.515 0.785 6.435 1.015 ;
        RECT 0.005 0.200 6.435 0.785 ;
        RECT 0.005 0.105 1.355 0.200 ;
        RECT 2.580 0.105 6.435 0.200 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.355 6.630 2.910 ;
        RECT -0.190 1.305 0.995 1.355 ;
        RECT 2.620 1.305 6.630 1.355 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 6.090 1.495 6.355 2.455 ;
        RECT 6.170 0.595 6.355 1.495 ;
        RECT 6.055 0.255 6.355 0.595 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.015 2.025 1.240 2.465 ;
        RECT 1.450 2.195 1.815 2.635 ;
        RECT 2.475 2.255 3.225 2.425 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.085 0.985 0.330 1.625 ;
        RECT 0.610 1.390 0.780 1.795 ;
        RECT 1.015 1.855 2.590 2.025 ;
        RECT 0.610 1.060 0.840 1.390 ;
        RECT 0.610 0.785 0.780 1.060 ;
        RECT 0.175 0.615 0.780 0.785 ;
        RECT 0.175 0.260 0.345 0.615 ;
        RECT 0.515 0.085 0.845 0.445 ;
        RECT 1.015 0.260 1.280 1.855 ;
        RECT 2.390 0.985 2.590 1.855 ;
        RECT 3.055 1.325 3.225 2.255 ;
        RECT 3.395 2.135 3.695 2.635 ;
        RECT 3.910 1.865 4.130 2.435 ;
        RECT 4.310 2.010 4.595 2.635 ;
        RECT 3.430 1.840 4.130 1.865 ;
        RECT 5.005 1.895 5.335 2.465 ;
        RECT 5.570 2.130 5.920 2.635 ;
        RECT 3.430 1.535 4.710 1.840 ;
        RECT 5.005 1.725 5.920 1.895 ;
        RECT 4.345 1.325 4.710 1.535 ;
        RECT 3.055 1.155 4.175 1.325 ;
        RECT 3.555 0.995 4.175 1.155 ;
        RECT 4.345 0.995 4.740 1.325 ;
        RECT 5.190 1.105 5.510 1.435 ;
        RECT 5.750 1.325 5.920 1.725 ;
        RECT 1.480 0.085 1.810 0.905 ;
        RECT 2.390 0.815 3.220 0.985 ;
        RECT 3.555 0.560 3.725 0.995 ;
        RECT 4.345 0.615 4.580 0.995 ;
        RECT 5.750 0.935 6.000 1.325 ;
        RECT 4.935 0.765 6.000 0.935 ;
        RECT 4.935 0.620 5.155 0.765 ;
        RECT 2.790 0.390 3.725 0.560 ;
        RECT 3.895 0.085 4.145 0.610 ;
        RECT 4.320 0.255 4.580 0.615 ;
        RECT 4.840 0.290 5.155 0.620 ;
        RECT 5.670 0.085 5.840 0.545 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 1.105 0.315 1.275 ;
        RECT 5.210 1.105 5.380 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
END sky130_fd_sc_hd__dlclkp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dlclkp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlclkp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER met1 ;
        RECT 0.090 1.260 0.380 1.305 ;
        RECT 5.150 1.260 5.440 1.305 ;
        RECT 0.090 1.120 5.440 1.260 ;
        RECT 0.090 1.075 0.380 1.120 ;
        RECT 5.150 1.075 5.440 1.120 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.530 1.435 2.215 1.685 ;
        RECT 1.985 0.285 2.215 1.435 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.395 0.880 2.440 1.145 ;
        RECT 3.680 0.880 4.655 1.015 ;
        RECT 1.395 0.785 4.655 0.880 ;
        RECT 5.515 0.785 6.895 1.015 ;
        RECT 0.005 0.200 6.895 0.785 ;
        RECT 0.005 0.105 1.355 0.200 ;
        RECT 2.585 0.105 6.895 0.200 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.355 7.090 2.910 ;
        RECT -0.190 1.305 0.995 1.355 ;
        RECT 2.625 1.305 7.090 1.355 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 6.095 1.495 6.360 2.455 ;
        RECT 6.165 0.595 6.360 1.495 ;
        RECT 6.060 0.255 6.360 0.595 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.015 2.025 1.240 2.465 ;
        RECT 1.455 2.195 1.820 2.635 ;
        RECT 2.480 2.255 3.230 2.425 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.090 0.985 0.330 1.625 ;
        RECT 0.610 1.390 0.780 1.795 ;
        RECT 1.015 1.855 2.645 2.025 ;
        RECT 0.610 1.060 0.840 1.390 ;
        RECT 0.610 0.785 0.780 1.060 ;
        RECT 0.175 0.615 0.780 0.785 ;
        RECT 0.175 0.260 0.345 0.615 ;
        RECT 0.515 0.085 0.845 0.445 ;
        RECT 1.015 0.260 1.280 1.855 ;
        RECT 2.395 0.985 2.645 1.855 ;
        RECT 3.060 1.325 3.230 2.255 ;
        RECT 3.400 2.135 3.700 2.635 ;
        RECT 3.915 1.865 4.135 2.435 ;
        RECT 4.315 2.010 4.600 2.635 ;
        RECT 3.435 1.840 4.135 1.865 ;
        RECT 5.010 1.895 5.340 2.465 ;
        RECT 5.575 2.130 5.925 2.635 ;
        RECT 3.435 1.535 4.735 1.840 ;
        RECT 5.010 1.725 5.925 1.895 ;
        RECT 3.060 1.155 4.180 1.325 ;
        RECT 3.555 0.995 4.180 1.155 ;
        RECT 4.350 0.995 4.735 1.535 ;
        RECT 5.210 1.105 5.485 1.435 ;
        RECT 5.755 1.325 5.925 1.725 ;
        RECT 6.530 1.485 6.810 2.635 ;
        RECT 1.485 0.085 1.815 0.905 ;
        RECT 2.395 0.815 3.225 0.985 ;
        RECT 3.555 0.560 3.725 0.995 ;
        RECT 4.350 0.615 4.585 0.995 ;
        RECT 5.755 0.935 5.995 1.325 ;
        RECT 4.930 0.765 5.995 0.935 ;
        RECT 4.930 0.620 5.150 0.765 ;
        RECT 2.795 0.390 3.725 0.560 ;
        RECT 3.895 0.085 4.145 0.610 ;
        RECT 4.315 0.255 4.585 0.615 ;
        RECT 4.835 0.290 5.150 0.620 ;
        RECT 5.675 0.085 5.845 0.545 ;
        RECT 6.530 0.085 6.810 0.885 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.150 1.105 0.320 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
  END
END sky130_fd_sc_hd__dlclkp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dlclkp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlclkp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.406500 ;
    PORT
      LAYER met1 ;
        RECT 0.090 1.260 0.380 1.305 ;
        RECT 5.170 1.260 5.460 1.305 ;
        RECT 0.090 1.120 5.460 1.260 ;
        RECT 0.090 1.075 0.380 1.120 ;
        RECT 5.170 1.075 5.460 1.120 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.530 0.765 1.950 1.015 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.750 0.785 7.810 1.015 ;
        RECT 0.005 0.105 7.810 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.039500 ;
    PORT
      LAYER li1 ;
        RECT 6.040 2.005 6.370 2.455 ;
        RECT 6.970 2.005 7.300 2.465 ;
        RECT 6.040 1.835 7.300 2.005 ;
        RECT 6.585 1.785 7.300 1.835 ;
        RECT 6.750 0.885 7.300 1.785 ;
        RECT 6.290 0.715 7.300 0.885 ;
        RECT 6.290 0.545 6.460 0.715 ;
        RECT 6.040 0.255 6.460 0.545 ;
        RECT 6.970 0.255 7.300 0.715 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.085 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.085 1.795 0.780 1.965 ;
        RECT 0.090 0.985 0.330 1.625 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.585 1.240 2.465 ;
        RECT 1.450 2.195 1.815 2.635 ;
        RECT 2.475 2.195 3.165 2.425 ;
        RECT 2.915 2.105 3.165 2.195 ;
        RECT 3.335 2.175 3.695 2.635 ;
        RECT 2.915 2.090 3.180 2.105 ;
        RECT 2.915 2.060 3.185 2.090 ;
        RECT 1.525 1.905 2.735 2.025 ;
        RECT 2.980 2.015 3.185 2.060 ;
        RECT 1.525 1.855 2.845 1.905 ;
        RECT 1.525 1.785 1.695 1.855 ;
        RECT 2.045 1.585 2.335 1.685 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 1.015 1.355 2.335 1.585 ;
        RECT 2.505 1.575 2.845 1.855 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.085 0.635 0.780 0.805 ;
        RECT 0.085 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.280 1.355 ;
        RECT 2.565 1.035 2.735 1.575 ;
        RECT 3.015 1.325 3.185 2.015 ;
        RECT 3.895 1.865 4.115 2.435 ;
        RECT 4.295 2.010 4.580 2.635 ;
        RECT 3.355 1.535 4.115 1.865 ;
        RECT 3.945 1.325 4.115 1.535 ;
        RECT 4.750 1.665 5.035 2.465 ;
        RECT 5.575 1.835 5.840 2.635 ;
        RECT 6.540 2.175 6.800 2.635 ;
        RECT 4.750 1.495 6.140 1.665 ;
        RECT 3.015 1.165 3.775 1.325 ;
        RECT 2.290 0.705 2.735 1.035 ;
        RECT 2.905 0.995 3.775 1.165 ;
        RECT 3.945 0.995 4.720 1.325 ;
        RECT 2.905 0.535 3.075 0.995 ;
        RECT 3.945 0.745 4.115 0.995 ;
        RECT 4.890 0.885 5.060 1.495 ;
        RECT 5.230 1.055 5.740 1.325 ;
        RECT 5.910 1.290 6.140 1.495 ;
        RECT 7.470 1.485 7.735 2.635 ;
        RECT 5.910 1.055 6.580 1.290 ;
        RECT 5.910 0.885 6.120 1.055 ;
        RECT 4.890 0.825 6.120 0.885 ;
        RECT 1.450 0.085 1.785 0.465 ;
        RECT 2.415 0.365 3.075 0.535 ;
        RECT 3.315 0.085 3.650 0.530 ;
        RECT 3.895 0.415 4.115 0.745 ;
        RECT 4.750 0.715 6.120 0.825 ;
        RECT 4.295 0.085 4.580 0.715 ;
        RECT 4.750 0.290 5.060 0.715 ;
        RECT 5.590 0.085 5.870 0.545 ;
        RECT 6.630 0.085 6.800 0.545 ;
        RECT 7.470 0.085 7.735 0.885 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.610 1.785 0.780 1.955 ;
        RECT 0.150 1.105 0.320 1.275 ;
        RECT 5.230 1.105 5.400 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
      LAYER met1 ;
        RECT 0.550 1.940 0.840 1.985 ;
        RECT 1.465 1.940 1.755 1.985 ;
        RECT 0.550 1.800 1.755 1.940 ;
        RECT 0.550 1.755 0.840 1.800 ;
        RECT 1.465 1.755 1.755 1.800 ;
  END
END sky130_fd_sc_hd__dlclkp_4

#--------EOF---------

MACRO sky130_fd_sc_hd__dlrbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.460 0.955 1.790 1.325 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 4.470 0.995 5.455 1.325 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.170 0.785 7.815 1.015 ;
        RECT 0.005 0.105 7.815 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 6.060 0.255 6.380 2.465 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 7.475 1.785 7.735 2.465 ;
        RECT 7.560 0.595 7.735 1.785 ;
        RECT 7.475 0.255 7.735 0.595 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.085 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.085 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.085 0.635 0.780 0.805 ;
        RECT 0.085 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.455 1.665 1.785 2.415 ;
        RECT 1.955 1.835 2.270 2.635 ;
        RECT 2.900 2.255 3.650 2.425 ;
        RECT 1.455 1.495 2.140 1.665 ;
        RECT 1.970 1.095 2.140 1.495 ;
        RECT 2.470 1.355 2.755 2.005 ;
        RECT 2.925 1.415 3.265 1.995 ;
        RECT 1.970 0.785 2.340 1.095 ;
        RECT 2.925 1.035 3.095 1.415 ;
        RECT 3.480 1.325 3.650 2.255 ;
        RECT 3.820 2.135 4.090 2.635 ;
        RECT 4.260 2.135 4.590 2.635 ;
        RECT 4.760 1.865 4.970 2.435 ;
        RECT 5.150 1.935 5.890 2.635 ;
        RECT 3.840 1.765 4.970 1.865 ;
        RECT 3.840 1.535 5.875 1.765 ;
        RECT 3.480 1.165 4.300 1.325 ;
        RECT 1.535 0.765 2.340 0.785 ;
        RECT 1.535 0.615 2.140 0.765 ;
        RECT 2.715 0.705 3.095 1.035 ;
        RECT 3.330 0.995 4.300 1.165 ;
        RECT 1.535 0.345 1.705 0.615 ;
        RECT 3.330 0.535 3.500 0.995 ;
        RECT 5.625 0.825 5.875 1.535 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 2.840 0.365 3.500 0.535 ;
        RECT 4.240 0.655 5.875 0.825 ;
        RECT 6.580 1.325 6.830 2.465 ;
        RECT 7.010 1.835 7.305 2.635 ;
        RECT 6.580 0.995 7.390 1.325 ;
        RECT 6.580 0.985 6.830 0.995 ;
        RECT 3.740 0.085 4.070 0.530 ;
        RECT 4.240 0.255 4.540 0.655 ;
        RECT 5.135 0.085 5.875 0.485 ;
        RECT 6.580 0.255 6.750 0.985 ;
        RECT 6.975 0.085 7.305 0.465 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.470 1.785 2.640 1.955 ;
        RECT 2.930 1.445 3.100 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.410 1.940 2.700 1.985 ;
        RECT 1.010 1.800 2.700 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.410 1.755 2.700 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.870 1.600 3.160 1.645 ;
        RECT 0.550 1.460 3.160 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.870 1.415 3.160 1.460 ;
  END
END sky130_fd_sc_hd__dlrbn_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dlrbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.460 0.955 1.790 1.325 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 4.390 0.995 5.140 1.325 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.170 0.785 8.265 1.015 ;
        RECT 0.005 0.105 8.265 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536250 ;
    PORT
      LAYER li1 ;
        RECT 5.650 1.660 5.915 2.465 ;
        RECT 5.650 1.495 5.975 1.660 ;
        RECT 5.790 1.325 5.975 1.495 ;
        RECT 5.790 0.885 6.355 1.325 ;
        RECT 5.790 0.860 5.975 0.885 ;
        RECT 5.740 0.825 5.975 0.860 ;
        RECT 5.650 0.685 5.975 0.825 ;
        RECT 5.650 0.655 5.950 0.685 ;
        RECT 5.650 0.415 5.910 0.655 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.453750 ;
    PORT
      LAYER li1 ;
        RECT 7.500 1.445 7.755 2.465 ;
        RECT 7.545 1.325 7.755 1.445 ;
        RECT 7.545 1.055 8.195 1.325 ;
        RECT 7.545 0.825 7.755 1.055 ;
        RECT 7.500 0.255 7.755 0.825 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.085 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.085 1.795 0.780 1.965 ;
        RECT 0.605 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.605 1.070 0.840 1.400 ;
        RECT 0.605 0.805 0.780 1.070 ;
        RECT 0.085 0.635 0.780 0.805 ;
        RECT 0.085 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.455 1.665 1.785 2.415 ;
        RECT 1.955 1.835 2.270 2.635 ;
        RECT 2.900 2.255 3.650 2.425 ;
        RECT 1.455 1.495 2.140 1.665 ;
        RECT 1.970 1.095 2.140 1.495 ;
        RECT 2.470 1.355 2.755 2.005 ;
        RECT 2.925 1.415 3.265 1.995 ;
        RECT 1.970 0.785 2.340 1.095 ;
        RECT 2.925 1.035 3.095 1.415 ;
        RECT 3.480 1.325 3.650 2.255 ;
        RECT 3.820 2.135 4.590 2.635 ;
        RECT 4.760 1.865 4.930 2.435 ;
        RECT 3.840 1.665 4.930 1.865 ;
        RECT 5.100 1.855 5.350 2.635 ;
        RECT 6.085 1.830 6.355 2.635 ;
        RECT 3.840 1.495 5.480 1.665 ;
        RECT 5.310 1.325 5.480 1.495 ;
        RECT 6.525 1.325 6.855 2.465 ;
        RECT 7.035 1.835 7.330 2.635 ;
        RECT 7.925 1.495 8.195 2.635 ;
        RECT 3.480 1.165 4.200 1.325 ;
        RECT 1.535 0.765 2.340 0.785 ;
        RECT 1.535 0.615 2.140 0.765 ;
        RECT 2.715 0.705 3.095 1.035 ;
        RECT 3.330 0.995 4.200 1.165 ;
        RECT 5.310 0.995 5.620 1.325 ;
        RECT 6.525 0.995 7.375 1.325 ;
        RECT 1.535 0.345 1.705 0.615 ;
        RECT 3.330 0.535 3.500 0.995 ;
        RECT 5.310 0.825 5.480 0.995 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 2.840 0.365 3.500 0.535 ;
        RECT 3.740 0.085 4.070 0.825 ;
        RECT 4.340 0.655 5.480 0.825 ;
        RECT 4.340 0.415 4.560 0.655 ;
        RECT 5.100 0.085 5.480 0.485 ;
        RECT 6.085 0.085 6.355 0.545 ;
        RECT 6.525 0.255 6.855 0.995 ;
        RECT 7.025 0.085 7.330 0.545 ;
        RECT 7.925 0.085 8.195 0.885 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.470 1.785 2.640 1.955 ;
        RECT 2.930 1.445 3.100 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.410 1.940 2.700 1.985 ;
        RECT 1.010 1.800 2.700 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.410 1.755 2.700 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.870 1.600 3.160 1.645 ;
        RECT 0.550 1.460 3.160 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.870 1.415 3.160 1.460 ;
  END
END sky130_fd_sc_hd__dlrbn_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dlrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.460 0.955 1.790 1.325 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.325 1.625 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 4.450 0.995 5.435 1.325 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.165 0.785 7.815 1.015 ;
        RECT 0.005 0.105 7.815 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 6.060 0.255 6.410 2.465 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 7.475 1.785 7.735 2.465 ;
        RECT 7.565 0.595 7.735 1.785 ;
        RECT 7.475 0.255 7.735 0.595 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.085 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.085 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.085 0.635 0.780 0.805 ;
        RECT 0.085 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.455 1.665 1.785 2.415 ;
        RECT 1.955 1.835 2.270 2.635 ;
        RECT 2.745 2.255 3.585 2.425 ;
        RECT 3.270 2.125 3.585 2.255 ;
        RECT 3.755 2.135 4.590 2.635 ;
        RECT 3.305 2.075 3.585 2.125 ;
        RECT 3.395 2.045 3.585 2.075 ;
        RECT 3.395 2.015 3.605 2.045 ;
        RECT 2.925 1.905 3.130 1.995 ;
        RECT 3.415 1.990 3.605 2.015 ;
        RECT 3.420 1.975 3.605 1.990 ;
        RECT 3.430 1.960 3.605 1.975 ;
        RECT 1.455 1.495 2.140 1.665 ;
        RECT 1.970 1.095 2.140 1.495 ;
        RECT 2.470 1.355 2.755 1.685 ;
        RECT 2.925 1.575 3.265 1.905 ;
        RECT 1.970 0.785 2.340 1.095 ;
        RECT 2.925 1.035 3.095 1.575 ;
        RECT 3.435 1.325 3.605 1.960 ;
        RECT 4.780 1.865 4.950 2.435 ;
        RECT 5.120 1.935 5.890 2.635 ;
        RECT 3.840 1.765 4.950 1.865 ;
        RECT 3.840 1.535 5.890 1.765 ;
        RECT 3.435 1.165 4.200 1.325 ;
        RECT 1.535 0.765 2.340 0.785 ;
        RECT 2.600 0.765 3.095 1.035 ;
        RECT 3.330 0.995 4.200 1.165 ;
        RECT 1.535 0.615 2.140 0.765 ;
        RECT 1.535 0.345 1.705 0.615 ;
        RECT 3.330 0.535 3.500 0.995 ;
        RECT 5.655 0.825 5.890 1.535 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 2.770 0.365 3.500 0.535 ;
        RECT 4.240 0.655 5.890 0.825 ;
        RECT 6.580 1.325 6.830 2.465 ;
        RECT 7.010 1.835 7.305 2.635 ;
        RECT 6.580 0.995 7.395 1.325 ;
        RECT 3.735 0.085 4.070 0.530 ;
        RECT 4.240 0.255 4.540 0.655 ;
        RECT 5.120 0.085 5.890 0.485 ;
        RECT 6.580 0.255 6.805 0.995 ;
        RECT 6.975 0.085 7.305 0.465 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.925 1.785 3.095 1.955 ;
        RECT 2.470 1.445 2.640 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.865 1.940 3.155 1.985 ;
        RECT 1.010 1.800 3.155 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.865 1.755 3.155 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.410 1.600 2.700 1.645 ;
        RECT 0.550 1.460 2.700 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.410 1.415 2.700 1.460 ;
  END
END sky130_fd_sc_hd__dlrbp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dlrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.460 0.955 1.790 1.325 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 4.400 0.995 5.150 1.325 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.170 0.785 8.275 1.015 ;
        RECT 0.005 0.105 8.275 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.478500 ;
    PORT
      LAYER li1 ;
        RECT 5.680 1.660 5.930 2.465 ;
        RECT 5.680 1.495 6.065 1.660 ;
        RECT 5.790 1.325 6.065 1.495 ;
        RECT 5.790 0.885 6.360 1.325 ;
        RECT 5.790 0.835 6.150 0.885 ;
        RECT 5.680 0.665 6.150 0.835 ;
        RECT 5.680 0.330 5.850 0.665 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 7.515 1.605 7.765 2.465 ;
        RECT 7.595 1.325 7.765 1.605 ;
        RECT 7.595 1.055 8.195 1.325 ;
        RECT 7.595 0.825 7.765 1.055 ;
        RECT 7.515 0.255 7.765 0.825 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.085 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.085 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.085 0.635 0.780 0.805 ;
        RECT 0.085 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.455 1.665 1.785 2.415 ;
        RECT 1.955 1.835 2.270 2.635 ;
        RECT 2.745 2.255 3.585 2.425 ;
        RECT 3.270 2.125 3.585 2.255 ;
        RECT 3.755 2.135 4.600 2.635 ;
        RECT 3.305 2.075 3.585 2.125 ;
        RECT 3.395 2.045 3.585 2.075 ;
        RECT 3.395 2.015 3.605 2.045 ;
        RECT 2.925 1.905 3.125 1.995 ;
        RECT 3.415 1.990 3.605 2.015 ;
        RECT 3.420 1.975 3.605 1.990 ;
        RECT 3.430 1.960 3.605 1.975 ;
        RECT 1.455 1.495 2.140 1.665 ;
        RECT 1.970 1.095 2.140 1.495 ;
        RECT 2.470 1.355 2.755 1.685 ;
        RECT 2.925 1.575 3.265 1.905 ;
        RECT 1.970 0.785 2.340 1.095 ;
        RECT 2.925 1.035 3.095 1.575 ;
        RECT 3.435 1.325 3.605 1.960 ;
        RECT 4.770 1.865 4.940 2.435 ;
        RECT 5.110 1.875 5.490 2.635 ;
        RECT 3.840 1.705 4.940 1.865 ;
        RECT 6.100 1.830 6.360 2.635 ;
        RECT 3.840 1.535 5.510 1.705 ;
        RECT 5.320 1.325 5.510 1.535 ;
        RECT 6.535 1.325 6.870 2.465 ;
        RECT 7.045 1.835 7.340 2.635 ;
        RECT 7.935 1.495 8.195 2.635 ;
        RECT 3.435 1.165 4.200 1.325 ;
        RECT 1.535 0.765 2.340 0.785 ;
        RECT 1.535 0.615 2.140 0.765 ;
        RECT 2.715 0.705 3.095 1.035 ;
        RECT 3.330 0.995 4.200 1.165 ;
        RECT 5.320 0.995 5.620 1.325 ;
        RECT 6.535 0.995 7.425 1.325 ;
        RECT 1.535 0.345 1.705 0.615 ;
        RECT 3.330 0.535 3.500 0.995 ;
        RECT 5.320 0.825 5.510 0.995 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 2.770 0.365 3.500 0.535 ;
        RECT 4.270 0.655 5.510 0.825 ;
        RECT 3.740 0.085 4.070 0.530 ;
        RECT 4.270 0.415 4.570 0.655 ;
        RECT 5.110 0.085 5.490 0.485 ;
        RECT 6.020 0.085 6.360 0.465 ;
        RECT 6.535 0.255 6.865 0.995 ;
        RECT 7.035 0.085 7.340 0.545 ;
        RECT 7.935 0.085 8.195 0.885 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.930 1.785 3.100 1.955 ;
        RECT 2.470 1.445 2.640 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.870 1.940 3.160 1.985 ;
        RECT 1.010 1.800 3.160 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.870 1.755 3.160 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.410 1.600 2.700 1.645 ;
        RECT 0.550 1.460 2.700 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.410 1.415 2.700 1.460 ;
  END
END sky130_fd_sc_hd__dlrbp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dlrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.460 0.955 1.790 1.325 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 4.500 0.995 5.435 1.325 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.170 0.785 6.435 1.015 ;
        RECT 0.005 0.105 6.435 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 6.095 0.415 6.355 2.455 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.175 0.635 0.780 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.455 1.665 1.785 2.415 ;
        RECT 1.955 1.835 2.270 2.635 ;
        RECT 2.900 2.255 3.650 2.425 ;
        RECT 1.455 1.495 2.140 1.665 ;
        RECT 1.970 1.095 2.140 1.495 ;
        RECT 2.470 1.355 2.755 2.005 ;
        RECT 2.925 1.415 3.265 1.995 ;
        RECT 1.970 0.785 2.340 1.095 ;
        RECT 2.925 1.035 3.095 1.415 ;
        RECT 3.480 1.325 3.650 2.255 ;
        RECT 3.820 2.135 4.110 2.635 ;
        RECT 4.300 2.135 4.580 2.635 ;
        RECT 4.750 1.865 4.940 2.465 ;
        RECT 5.110 2.135 5.925 2.635 ;
        RECT 3.820 1.535 5.925 1.865 ;
        RECT 3.480 1.245 4.330 1.325 ;
        RECT 1.535 0.765 2.340 0.785 ;
        RECT 1.535 0.615 2.140 0.765 ;
        RECT 2.715 0.705 3.095 1.035 ;
        RECT 3.330 1.025 4.330 1.245 ;
        RECT 1.535 0.345 1.705 0.615 ;
        RECT 3.330 0.535 3.500 1.025 ;
        RECT 5.605 0.825 5.925 1.535 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 2.840 0.365 3.500 0.535 ;
        RECT 4.240 0.655 5.925 0.825 ;
        RECT 3.740 0.085 4.070 0.530 ;
        RECT 4.240 0.255 4.590 0.655 ;
        RECT 5.095 0.085 5.925 0.485 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.470 1.785 2.640 1.955 ;
        RECT 2.930 1.445 3.100 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.410 1.940 2.700 1.985 ;
        RECT 1.010 1.800 2.700 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.410 1.755 2.700 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.870 1.600 3.160 1.645 ;
        RECT 0.550 1.460 3.160 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.870 1.415 3.160 1.460 ;
  END
END sky130_fd_sc_hd__dlrtn_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dlrtn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.460 0.955 1.790 1.325 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 4.480 0.995 5.170 1.325 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.165 0.785 6.435 1.015 ;
        RECT 0.005 0.105 6.435 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.480500 ;
    PORT
      LAYER li1 ;
        RECT 5.655 1.875 5.925 2.465 ;
        RECT 5.755 1.500 5.925 1.875 ;
        RECT 5.755 1.425 6.355 1.500 ;
        RECT 5.760 1.415 6.355 1.425 ;
        RECT 5.765 1.410 6.355 1.415 ;
        RECT 5.775 1.385 6.355 1.410 ;
        RECT 5.785 0.890 6.355 1.385 ;
        RECT 5.770 0.865 6.355 0.890 ;
        RECT 5.755 0.765 6.355 0.865 ;
        RECT 5.755 0.485 5.925 0.765 ;
        RECT 5.595 0.255 5.925 0.485 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.175 0.635 0.780 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.455 1.665 1.785 2.415 ;
        RECT 1.955 1.835 2.270 2.635 ;
        RECT 2.775 2.255 3.605 2.425 ;
        RECT 1.455 1.495 2.140 1.665 ;
        RECT 1.960 1.095 2.140 1.495 ;
        RECT 2.470 1.355 2.755 2.005 ;
        RECT 2.925 1.415 3.265 1.995 ;
        RECT 2.925 1.145 3.095 1.415 ;
        RECT 3.435 1.325 3.605 2.255 ;
        RECT 3.800 2.135 4.110 2.635 ;
        RECT 4.280 2.135 4.560 2.635 ;
        RECT 4.730 1.865 4.920 2.465 ;
        RECT 5.090 1.875 5.460 2.635 ;
        RECT 3.820 1.705 4.920 1.865 ;
        RECT 3.820 1.535 5.585 1.705 ;
        RECT 6.095 1.670 6.355 2.635 ;
        RECT 5.415 1.325 5.585 1.535 ;
        RECT 3.435 1.245 4.310 1.325 ;
        RECT 1.960 0.785 2.340 1.095 ;
        RECT 1.535 0.765 2.340 0.785 ;
        RECT 1.535 0.615 2.140 0.765 ;
        RECT 2.675 0.705 3.095 1.145 ;
        RECT 3.330 1.025 4.310 1.245 ;
        RECT 1.535 0.345 1.705 0.615 ;
        RECT 3.330 0.535 3.500 1.025 ;
        RECT 5.350 0.995 5.615 1.325 ;
        RECT 5.415 0.825 5.585 0.995 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 2.810 0.365 3.500 0.535 ;
        RECT 4.240 0.655 5.585 0.825 ;
        RECT 3.735 0.085 4.070 0.530 ;
        RECT 4.240 0.255 4.590 0.655 ;
        RECT 5.095 0.085 5.425 0.485 ;
        RECT 6.095 0.085 6.355 0.595 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.470 1.785 2.640 1.955 ;
        RECT 2.930 1.445 3.100 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.410 1.940 2.700 1.985 ;
        RECT 1.010 1.800 2.700 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.410 1.755 2.700 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.870 1.600 3.160 1.645 ;
        RECT 0.550 1.460 3.160 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.870 1.415 3.160 1.460 ;
  END
END sky130_fd_sc_hd__dlrtn_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dlrtn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.465 0.955 1.795 1.325 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE_N
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 4.505 0.995 5.145 1.325 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.175 0.785 7.355 1.015 ;
        RECT 0.005 0.105 7.355 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.014750 ;
    PORT
      LAYER li1 ;
        RECT 5.680 1.875 5.965 2.465 ;
        RECT 5.795 1.325 5.965 1.875 ;
        RECT 6.575 1.325 6.775 2.465 ;
        RECT 5.795 0.765 7.275 1.325 ;
        RECT 5.795 0.485 5.965 0.765 ;
        RECT 5.610 0.255 5.965 0.485 ;
        RECT 6.575 0.255 6.775 0.765 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.175 0.635 0.780 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.460 1.665 1.790 2.415 ;
        RECT 1.960 1.835 2.275 2.635 ;
        RECT 2.905 2.255 3.655 2.425 ;
        RECT 1.460 1.495 2.145 1.665 ;
        RECT 1.975 1.095 2.145 1.495 ;
        RECT 2.475 1.355 2.760 2.005 ;
        RECT 2.930 1.415 3.270 1.995 ;
        RECT 1.975 0.785 2.345 1.095 ;
        RECT 2.930 1.035 3.100 1.415 ;
        RECT 3.485 1.325 3.655 2.255 ;
        RECT 3.825 2.135 4.115 2.635 ;
        RECT 4.305 2.135 4.585 2.635 ;
        RECT 4.755 1.865 4.945 2.465 ;
        RECT 5.115 1.875 5.485 2.635 ;
        RECT 3.825 1.705 4.945 1.865 ;
        RECT 3.825 1.535 5.625 1.705 ;
        RECT 3.485 1.245 4.315 1.325 ;
        RECT 1.540 0.765 2.345 0.785 ;
        RECT 1.540 0.615 2.145 0.765 ;
        RECT 2.720 0.705 3.100 1.035 ;
        RECT 3.335 1.025 4.315 1.245 ;
        RECT 1.540 0.345 1.710 0.615 ;
        RECT 3.335 0.535 3.505 1.025 ;
        RECT 5.455 0.825 5.625 1.535 ;
        RECT 6.135 1.495 6.405 2.635 ;
        RECT 6.945 1.495 7.275 2.635 ;
        RECT 1.880 0.085 2.210 0.445 ;
        RECT 2.845 0.365 3.505 0.535 ;
        RECT 4.245 0.655 5.625 0.825 ;
        RECT 3.745 0.085 4.075 0.530 ;
        RECT 4.245 0.255 4.595 0.655 ;
        RECT 5.100 0.085 5.440 0.485 ;
        RECT 6.135 0.085 6.405 0.595 ;
        RECT 6.945 0.085 7.275 0.595 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.475 1.785 2.645 1.955 ;
        RECT 2.935 1.445 3.105 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.415 1.940 2.705 1.985 ;
        RECT 1.010 1.800 2.705 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.415 1.755 2.705 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.875 1.600 3.165 1.645 ;
        RECT 0.550 1.460 3.165 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.875 1.415 3.165 1.460 ;
  END
END sky130_fd_sc_hd__dlrtn_4

#--------EOF---------

MACRO sky130_fd_sc_hd__dlrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.435 0.955 1.765 1.325 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.325 1.625 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 4.745 0.995 5.075 1.325 ;
        RECT 4.745 0.345 4.975 0.995 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.105 0.785 5.975 1.015 ;
        RECT 0.005 0.105 5.975 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 5.635 1.670 5.895 2.455 ;
        RECT 5.725 0.745 5.895 1.670 ;
        RECT 5.610 0.345 5.895 0.745 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.085 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.085 1.795 0.775 1.965 ;
        RECT 0.605 1.400 0.775 1.795 ;
        RECT 1.015 1.685 1.235 2.465 ;
        RECT 0.605 1.070 0.835 1.400 ;
        RECT 0.605 0.805 0.775 1.070 ;
        RECT 0.170 0.635 0.775 0.805 ;
        RECT 0.170 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.430 1.665 1.785 2.415 ;
        RECT 1.955 1.835 2.245 2.635 ;
        RECT 2.810 2.255 3.625 2.425 ;
        RECT 2.900 1.785 3.265 1.995 ;
        RECT 1.430 1.495 2.115 1.665 ;
        RECT 1.945 1.095 2.115 1.495 ;
        RECT 2.445 1.625 2.760 1.685 ;
        RECT 3.005 1.635 3.265 1.785 ;
        RECT 2.445 1.355 2.835 1.625 ;
        RECT 3.005 1.095 3.245 1.635 ;
        RECT 3.455 1.325 3.625 2.255 ;
        RECT 3.930 2.135 4.445 2.635 ;
        RECT 4.625 1.865 4.965 2.435 ;
        RECT 5.135 1.915 5.465 2.635 ;
        RECT 3.815 1.735 4.965 1.865 ;
        RECT 3.815 1.535 5.465 1.735 ;
        RECT 4.345 1.505 5.465 1.535 ;
        RECT 3.455 1.165 4.175 1.325 ;
        RECT 1.945 0.785 2.335 1.095 ;
        RECT 1.510 0.765 2.335 0.785 ;
        RECT 2.690 0.765 3.245 1.095 ;
        RECT 3.415 0.995 4.175 1.165 ;
        RECT 1.510 0.615 2.115 0.765 ;
        RECT 1.510 0.345 1.705 0.615 ;
        RECT 3.415 0.535 3.585 0.995 ;
        RECT 4.345 0.805 4.575 1.505 ;
        RECT 5.245 1.325 5.465 1.505 ;
        RECT 5.245 0.995 5.555 1.325 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 2.815 0.365 3.585 0.535 ;
        RECT 3.755 0.085 4.025 0.610 ;
        RECT 4.195 0.295 4.575 0.805 ;
        RECT 5.155 0.085 5.440 0.715 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.605 1.445 0.775 1.615 ;
        RECT 1.065 1.785 1.235 1.955 ;
        RECT 2.925 1.785 3.095 1.955 ;
        RECT 2.445 1.445 2.615 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
      LAYER met1 ;
        RECT 1.005 1.940 1.295 1.985 ;
        RECT 2.865 1.940 3.155 1.985 ;
        RECT 1.005 1.800 3.155 1.940 ;
        RECT 1.005 1.755 1.295 1.800 ;
        RECT 2.865 1.755 3.155 1.800 ;
        RECT 0.545 1.600 0.835 1.645 ;
        RECT 2.385 1.600 2.675 1.645 ;
        RECT 0.545 1.460 2.675 1.600 ;
        RECT 0.545 1.415 0.835 1.460 ;
        RECT 2.385 1.415 2.675 1.460 ;
  END
END sky130_fd_sc_hd__dlrtp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dlrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.440 0.955 1.770 1.325 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.985 0.330 1.625 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 4.480 1.035 5.240 1.325 ;
        RECT 4.480 0.995 4.815 1.035 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.160 0.785 6.435 1.015 ;
        RECT 0.005 0.105 6.435 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.480500 ;
    PORT
      LAYER li1 ;
        RECT 5.655 1.875 5.925 2.465 ;
        RECT 5.755 1.500 5.925 1.875 ;
        RECT 5.755 1.425 6.355 1.500 ;
        RECT 5.760 1.415 6.355 1.425 ;
        RECT 5.765 1.410 6.355 1.415 ;
        RECT 5.775 1.385 6.355 1.410 ;
        RECT 5.785 0.890 6.355 1.385 ;
        RECT 5.770 0.865 6.355 0.890 ;
        RECT 5.755 0.765 6.355 0.865 ;
        RECT 5.755 0.485 5.925 0.765 ;
        RECT 5.595 0.255 5.925 0.485 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.085 0.635 0.780 0.805 ;
        RECT 0.085 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.435 1.665 1.785 2.415 ;
        RECT 1.955 1.835 2.250 2.635 ;
        RECT 2.770 2.255 3.580 2.425 ;
        RECT 3.410 2.085 3.580 2.255 ;
        RECT 3.750 2.175 4.090 2.635 ;
        RECT 4.280 2.135 4.560 2.635 ;
        RECT 3.410 2.000 3.605 2.085 ;
        RECT 3.415 1.995 3.605 2.000 ;
        RECT 2.905 1.910 3.175 1.995 ;
        RECT 3.420 1.985 3.605 1.995 ;
        RECT 2.905 1.780 3.265 1.910 ;
        RECT 1.435 1.495 2.120 1.665 ;
        RECT 1.950 1.095 2.120 1.495 ;
        RECT 2.450 1.355 2.755 1.685 ;
        RECT 2.930 1.570 3.265 1.780 ;
        RECT 1.950 0.785 2.335 1.095 ;
        RECT 2.930 1.040 3.100 1.570 ;
        RECT 3.435 1.325 3.605 1.985 ;
        RECT 4.800 1.865 4.970 2.465 ;
        RECT 5.140 1.875 5.485 2.635 ;
        RECT 3.775 1.705 4.970 1.865 ;
        RECT 3.775 1.535 5.585 1.705 ;
        RECT 6.095 1.670 6.355 2.635 ;
        RECT 5.415 1.325 5.585 1.535 ;
        RECT 1.515 0.765 2.335 0.785 ;
        RECT 1.515 0.615 2.120 0.765 ;
        RECT 2.585 0.735 3.100 1.040 ;
        RECT 3.270 0.995 4.220 1.325 ;
        RECT 5.415 0.995 5.615 1.325 ;
        RECT 1.515 0.345 1.705 0.615 ;
        RECT 3.270 0.535 3.445 0.995 ;
        RECT 5.415 0.865 5.585 0.995 ;
        RECT 4.955 0.825 5.585 0.865 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 2.770 0.365 3.445 0.535 ;
        RECT 4.240 0.695 5.585 0.825 ;
        RECT 4.240 0.655 5.095 0.695 ;
        RECT 3.720 0.085 4.060 0.530 ;
        RECT 4.240 0.255 4.580 0.655 ;
        RECT 5.255 0.085 5.425 0.525 ;
        RECT 6.095 0.085 6.355 0.595 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.925 1.785 3.095 1.955 ;
        RECT 2.450 1.445 2.620 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.865 1.940 3.155 1.985 ;
        RECT 1.010 1.800 3.155 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.865 1.755 3.155 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.390 1.600 2.680 1.645 ;
        RECT 0.550 1.460 2.680 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.390 1.415 2.680 1.460 ;
  END
END sky130_fd_sc_hd__dlrtp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dlrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlrtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.465 0.955 1.795 1.325 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 4.505 0.995 5.145 1.325 ;
    END
  END RESET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.175 0.785 7.355 1.015 ;
        RECT 0.005 0.105 7.355 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.014750 ;
    PORT
      LAYER li1 ;
        RECT 5.680 1.875 5.965 2.465 ;
        RECT 5.795 1.325 5.965 1.875 ;
        RECT 6.575 1.325 6.775 2.465 ;
        RECT 5.795 0.765 7.275 1.325 ;
        RECT 5.795 0.485 5.965 0.765 ;
        RECT 5.610 0.255 5.965 0.485 ;
        RECT 6.575 0.255 6.775 0.765 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.175 0.635 0.780 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.460 1.665 1.790 2.415 ;
        RECT 1.960 1.835 2.275 2.635 ;
        RECT 2.905 2.255 3.655 2.425 ;
        RECT 1.460 1.495 2.145 1.665 ;
        RECT 1.975 1.095 2.145 1.495 ;
        RECT 2.475 1.355 2.760 1.685 ;
        RECT 2.930 1.575 3.270 1.995 ;
        RECT 1.975 0.785 2.345 1.095 ;
        RECT 2.930 1.035 3.100 1.575 ;
        RECT 3.485 1.325 3.655 2.255 ;
        RECT 3.825 2.135 4.115 2.635 ;
        RECT 4.305 2.135 4.585 2.635 ;
        RECT 4.755 1.865 4.945 2.465 ;
        RECT 5.115 1.875 5.485 2.635 ;
        RECT 3.825 1.705 4.945 1.865 ;
        RECT 3.825 1.535 5.625 1.705 ;
        RECT 3.485 1.165 4.235 1.325 ;
        RECT 1.540 0.765 2.345 0.785 ;
        RECT 1.540 0.615 2.145 0.765 ;
        RECT 2.720 0.705 3.100 1.035 ;
        RECT 3.335 0.995 4.235 1.165 ;
        RECT 1.540 0.345 1.710 0.615 ;
        RECT 3.335 0.535 3.505 0.995 ;
        RECT 5.455 0.825 5.625 1.535 ;
        RECT 6.135 1.495 6.405 2.635 ;
        RECT 6.945 1.495 7.275 2.635 ;
        RECT 1.880 0.085 2.210 0.445 ;
        RECT 2.845 0.365 3.505 0.535 ;
        RECT 4.265 0.655 5.625 0.825 ;
        RECT 3.745 0.085 4.075 0.530 ;
        RECT 4.265 0.255 4.595 0.655 ;
        RECT 5.100 0.085 5.440 0.485 ;
        RECT 6.135 0.085 6.405 0.595 ;
        RECT 6.945 0.085 7.275 0.595 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.935 1.785 3.105 1.955 ;
        RECT 2.475 1.445 2.645 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.875 1.940 3.165 1.985 ;
        RECT 1.010 1.800 3.165 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.875 1.755 3.165 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.415 1.600 2.705 1.645 ;
        RECT 0.550 1.460 2.705 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.415 1.415 2.705 1.460 ;
  END
END sky130_fd_sc_hd__dlrtp_4

#--------EOF---------

MACRO sky130_fd_sc_hd__dlxbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxbn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.445 0.955 1.785 1.325 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.985 0.330 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.130 0.785 6.895 1.015 ;
        RECT 0.005 0.105 6.895 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 5.140 1.670 5.480 2.465 ;
        RECT 5.310 0.745 5.480 1.670 ;
        RECT 5.140 0.415 5.480 0.745 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 6.555 1.505 6.815 2.465 ;
        RECT 6.625 0.825 6.815 1.505 ;
        RECT 6.555 0.255 6.815 0.825 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.175 0.635 0.780 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.480 1.665 1.810 2.415 ;
        RECT 1.980 1.835 2.295 2.635 ;
        RECT 2.920 2.130 3.610 2.275 ;
        RECT 3.780 2.175 3.950 2.635 ;
        RECT 2.920 2.115 3.615 2.130 ;
        RECT 2.920 2.105 3.620 2.115 ;
        RECT 3.360 2.090 3.625 2.105 ;
        RECT 3.360 2.075 3.630 2.090 ;
        RECT 3.375 2.060 3.630 2.075 ;
        RECT 3.420 2.030 3.630 2.060 ;
        RECT 3.430 2.015 3.630 2.030 ;
        RECT 1.480 1.495 2.165 1.665 ;
        RECT 1.995 1.235 2.165 1.495 ;
        RECT 2.495 1.355 2.780 2.005 ;
        RECT 2.950 1.415 3.290 1.910 ;
        RECT 1.995 0.905 2.365 1.235 ;
        RECT 2.950 1.035 3.120 1.415 ;
        RECT 3.460 1.325 3.630 2.015 ;
        RECT 4.300 1.865 4.550 2.435 ;
        RECT 3.800 1.620 4.550 1.865 ;
        RECT 4.720 1.830 4.970 2.635 ;
        RECT 3.800 1.535 4.580 1.620 ;
        RECT 4.395 1.325 4.580 1.535 ;
        RECT 5.660 1.325 5.910 2.465 ;
        RECT 6.090 1.835 6.385 2.635 ;
        RECT 3.460 1.165 4.225 1.325 ;
        RECT 1.995 0.785 2.165 0.905 ;
        RECT 1.535 0.615 2.165 0.785 ;
        RECT 2.565 0.705 3.120 1.035 ;
        RECT 3.355 0.995 4.225 1.165 ;
        RECT 4.395 0.995 5.140 1.325 ;
        RECT 5.660 0.995 6.455 1.325 ;
        RECT 1.535 0.345 1.705 0.615 ;
        RECT 3.355 0.535 3.525 0.995 ;
        RECT 4.395 0.840 4.580 0.995 ;
        RECT 4.300 0.660 4.580 0.840 ;
        RECT 1.875 0.085 2.230 0.445 ;
        RECT 2.790 0.365 3.525 0.535 ;
        RECT 3.765 0.085 4.095 0.610 ;
        RECT 4.300 0.415 4.470 0.660 ;
        RECT 4.640 0.085 4.970 0.495 ;
        RECT 5.660 0.255 5.910 0.995 ;
        RECT 6.090 0.085 6.385 0.545 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.495 1.785 2.665 1.955 ;
        RECT 2.955 1.445 3.125 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.435 1.940 2.725 1.985 ;
        RECT 1.010 1.800 2.725 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.435 1.755 2.725 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.895 1.600 3.185 1.645 ;
        RECT 0.550 1.460 3.185 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.895 1.415 3.185 1.460 ;
  END
END sky130_fd_sc_hd__dlxbn_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dlxbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxbn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.480 0.955 1.810 1.325 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.190 0.785 7.815 1.015 ;
        RECT 0.005 0.105 7.815 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 5.215 1.710 5.465 2.455 ;
        RECT 5.215 1.495 5.500 1.710 ;
        RECT 5.330 1.325 5.500 1.495 ;
        RECT 5.330 0.995 5.905 1.325 ;
        RECT 5.330 0.825 5.500 0.995 ;
        RECT 5.215 0.660 5.500 0.825 ;
        RECT 5.215 0.415 5.465 0.660 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.453750 ;
    PORT
      LAYER li1 ;
        RECT 7.050 1.445 7.305 2.465 ;
        RECT 7.095 1.325 7.305 1.445 ;
        RECT 7.095 1.055 7.735 1.325 ;
        RECT 7.095 0.825 7.305 1.055 ;
        RECT 7.050 0.255 7.305 0.825 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.175 0.635 0.780 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.475 1.665 1.805 2.415 ;
        RECT 1.975 1.835 2.290 2.635 ;
        RECT 2.920 2.255 3.670 2.425 ;
        RECT 1.475 1.495 2.160 1.665 ;
        RECT 1.990 1.095 2.160 1.495 ;
        RECT 2.490 1.355 2.775 2.005 ;
        RECT 2.945 1.415 3.285 1.995 ;
        RECT 1.990 0.785 2.360 1.095 ;
        RECT 2.945 1.035 3.115 1.415 ;
        RECT 3.500 1.325 3.670 2.255 ;
        RECT 3.840 2.135 4.140 2.635 ;
        RECT 4.360 1.865 4.580 2.435 ;
        RECT 3.860 1.535 4.580 1.865 ;
        RECT 4.410 1.325 4.580 1.535 ;
        RECT 4.760 1.495 5.045 2.635 ;
        RECT 5.635 1.835 5.905 2.635 ;
        RECT 6.075 1.325 6.405 2.465 ;
        RECT 6.585 1.835 6.880 2.635 ;
        RECT 7.475 1.495 7.735 2.635 ;
        RECT 3.500 1.165 4.220 1.325 ;
        RECT 1.555 0.765 2.360 0.785 ;
        RECT 1.555 0.615 2.160 0.765 ;
        RECT 2.735 0.705 3.115 1.035 ;
        RECT 3.350 0.995 4.220 1.165 ;
        RECT 4.410 0.995 5.160 1.325 ;
        RECT 6.075 0.995 6.925 1.325 ;
        RECT 1.555 0.345 1.725 0.615 ;
        RECT 3.350 0.535 3.520 0.995 ;
        RECT 4.410 0.825 4.580 0.995 ;
        RECT 1.895 0.085 2.225 0.445 ;
        RECT 2.860 0.365 3.520 0.535 ;
        RECT 3.760 0.085 4.090 0.825 ;
        RECT 4.360 0.415 4.580 0.825 ;
        RECT 4.760 0.085 5.045 0.825 ;
        RECT 5.635 0.085 5.905 0.545 ;
        RECT 6.075 0.255 6.405 0.995 ;
        RECT 6.585 0.085 6.880 0.545 ;
        RECT 7.475 0.085 7.735 0.885 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.490 1.785 2.660 1.955 ;
        RECT 2.950 1.445 3.120 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.430 1.940 2.720 1.985 ;
        RECT 1.010 1.800 2.720 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.430 1.755 2.720 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.890 1.600 3.180 1.645 ;
        RECT 0.550 1.460 3.180 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.890 1.415 3.180 1.460 ;
  END
END sky130_fd_sc_hd__dlxbn_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dlxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.355 0.955 1.685 1.325 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.130 0.785 6.895 1.015 ;
        RECT 0.005 0.105 6.895 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 5.140 1.670 5.490 2.455 ;
        RECT 5.320 0.820 5.490 1.670 ;
        RECT 5.140 0.255 5.490 0.820 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 6.555 1.445 6.815 2.465 ;
        RECT 6.600 0.825 6.815 1.445 ;
        RECT 6.555 0.255 6.815 0.825 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.175 0.635 0.780 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.430 1.665 1.795 2.415 ;
        RECT 1.965 1.835 2.245 2.635 ;
        RECT 2.750 2.255 3.610 2.425 ;
        RECT 3.425 2.090 3.610 2.255 ;
        RECT 3.780 2.175 3.980 2.635 ;
        RECT 3.425 2.065 3.630 2.090 ;
        RECT 3.425 2.035 3.650 2.065 ;
        RECT 3.430 2.020 3.650 2.035 ;
        RECT 3.435 2.010 3.650 2.020 ;
        RECT 3.440 1.995 3.650 2.010 ;
        RECT 2.965 1.910 3.195 1.995 ;
        RECT 1.430 1.495 2.115 1.665 ;
        RECT 1.855 1.235 2.115 1.495 ;
        RECT 2.465 1.355 2.795 1.685 ;
        RECT 2.965 1.575 3.290 1.910 ;
        RECT 1.855 0.875 2.335 1.235 ;
        RECT 2.965 1.065 3.135 1.575 ;
        RECT 3.460 1.325 3.650 1.995 ;
        RECT 4.285 1.865 4.515 2.435 ;
        RECT 3.820 1.535 4.515 1.865 ;
        RECT 4.685 1.570 4.970 2.635 ;
        RECT 4.345 1.325 4.515 1.535 ;
        RECT 5.660 1.325 5.910 2.465 ;
        RECT 6.090 1.835 6.385 2.635 ;
        RECT 3.460 1.165 4.175 1.325 ;
        RECT 1.855 0.785 2.135 0.875 ;
        RECT 1.510 0.615 2.135 0.785 ;
        RECT 2.580 0.705 3.135 1.065 ;
        RECT 3.305 0.995 4.175 1.165 ;
        RECT 4.345 0.995 5.150 1.325 ;
        RECT 5.660 0.995 6.430 1.325 ;
        RECT 1.510 0.345 1.705 0.615 ;
        RECT 3.305 0.535 3.475 0.995 ;
        RECT 4.345 0.745 4.550 0.995 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 2.800 0.365 3.475 0.535 ;
        RECT 3.700 0.085 4.045 0.530 ;
        RECT 4.285 0.415 4.550 0.745 ;
        RECT 4.720 0.085 4.970 0.715 ;
        RECT 5.660 0.255 5.910 0.995 ;
        RECT 6.090 0.085 6.385 0.545 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.965 1.785 3.135 1.955 ;
        RECT 2.555 1.445 2.725 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.905 1.940 3.195 1.985 ;
        RECT 1.010 1.800 3.195 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.905 1.755 3.195 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.495 1.600 2.785 1.645 ;
        RECT 0.550 1.460 2.785 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.495 1.415 2.785 1.460 ;
  END
END sky130_fd_sc_hd__dlxbp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dlxtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.435 0.955 1.765 1.325 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.125 0.785 5.515 1.015 ;
        RECT 0.005 0.105 5.515 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 5.175 1.670 5.435 2.455 ;
        RECT 5.265 0.745 5.435 1.670 ;
        RECT 5.175 0.415 5.435 0.745 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.175 0.635 0.780 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.430 1.665 1.785 2.415 ;
        RECT 1.955 1.835 2.245 2.635 ;
        RECT 2.745 2.255 3.605 2.425 ;
        RECT 3.295 2.105 3.605 2.255 ;
        RECT 3.775 2.175 4.095 2.635 ;
        RECT 3.295 2.090 3.620 2.105 ;
        RECT 3.390 2.085 3.620 2.090 ;
        RECT 3.390 2.065 3.630 2.085 ;
        RECT 3.390 2.045 3.645 2.065 ;
        RECT 3.405 2.035 3.645 2.045 ;
        RECT 3.430 2.010 3.645 2.035 ;
        RECT 1.430 1.495 2.115 1.665 ;
        RECT 1.945 1.235 2.115 1.495 ;
        RECT 2.445 1.355 2.780 2.005 ;
        RECT 2.950 1.560 3.285 1.910 ;
        RECT 1.945 0.785 2.320 1.235 ;
        RECT 2.950 1.040 3.265 1.560 ;
        RECT 3.455 1.450 3.645 2.010 ;
        RECT 4.295 1.865 4.540 2.435 ;
        RECT 3.815 1.535 4.540 1.865 ;
        RECT 4.720 1.570 5.005 2.635 ;
        RECT 1.510 0.765 2.320 0.785 ;
        RECT 1.510 0.615 2.115 0.765 ;
        RECT 2.560 0.735 3.265 1.040 ;
        RECT 3.435 1.325 3.645 1.450 ;
        RECT 4.370 1.325 4.540 1.535 ;
        RECT 3.435 0.995 4.200 1.325 ;
        RECT 4.370 0.995 5.095 1.325 ;
        RECT 1.510 0.345 1.705 0.615 ;
        RECT 3.435 0.535 3.605 0.995 ;
        RECT 4.370 0.720 4.540 0.995 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 2.765 0.365 3.605 0.535 ;
        RECT 3.775 0.085 4.045 0.545 ;
        RECT 4.295 0.260 4.540 0.720 ;
        RECT 4.755 0.085 4.980 0.715 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.445 1.785 2.615 1.955 ;
        RECT 2.950 1.445 3.120 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.385 1.940 2.675 1.985 ;
        RECT 1.010 1.800 2.675 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.385 1.755 2.675 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.890 1.600 3.180 1.645 ;
        RECT 0.550 1.460 3.180 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.890 1.415 3.180 1.460 ;
  END
END sky130_fd_sc_hd__dlxtn_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dlxtn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.480 0.955 1.810 1.325 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.190 0.785 5.975 1.015 ;
        RECT 0.005 0.105 5.975 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 5.215 1.640 5.465 2.455 ;
        RECT 5.215 1.495 5.500 1.640 ;
        RECT 5.330 1.325 5.500 1.495 ;
        RECT 5.330 0.995 5.895 1.325 ;
        RECT 5.330 0.825 5.500 0.995 ;
        RECT 5.215 0.685 5.500 0.825 ;
        RECT 5.215 0.415 5.465 0.685 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.175 0.635 0.780 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.475 1.665 1.805 2.415 ;
        RECT 1.975 1.835 2.290 2.635 ;
        RECT 2.920 2.255 3.670 2.425 ;
        RECT 1.475 1.495 2.160 1.665 ;
        RECT 1.990 1.095 2.160 1.495 ;
        RECT 2.490 1.355 2.775 2.005 ;
        RECT 2.945 1.415 3.285 1.995 ;
        RECT 1.990 0.785 2.360 1.095 ;
        RECT 2.945 1.035 3.115 1.415 ;
        RECT 3.500 1.325 3.670 2.255 ;
        RECT 3.840 2.135 4.140 2.635 ;
        RECT 4.360 1.865 4.580 2.435 ;
        RECT 3.860 1.535 4.580 1.865 ;
        RECT 4.410 1.325 4.580 1.535 ;
        RECT 4.760 1.495 5.045 2.635 ;
        RECT 5.635 1.755 5.895 2.635 ;
        RECT 3.500 1.165 4.220 1.325 ;
        RECT 1.555 0.765 2.360 0.785 ;
        RECT 1.555 0.615 2.160 0.765 ;
        RECT 2.735 0.705 3.115 1.035 ;
        RECT 3.350 0.995 4.220 1.165 ;
        RECT 4.410 0.995 5.160 1.325 ;
        RECT 1.555 0.345 1.725 0.615 ;
        RECT 3.350 0.535 3.520 0.995 ;
        RECT 4.410 0.825 4.580 0.995 ;
        RECT 1.895 0.085 2.225 0.445 ;
        RECT 2.860 0.365 3.520 0.535 ;
        RECT 3.760 0.085 4.090 0.825 ;
        RECT 4.360 0.415 4.580 0.825 ;
        RECT 4.760 0.085 5.045 0.825 ;
        RECT 5.635 0.085 5.895 0.550 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.490 1.785 2.660 1.955 ;
        RECT 2.950 1.445 3.120 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.430 1.940 2.720 1.985 ;
        RECT 1.010 1.800 2.720 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.430 1.755 2.720 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.890 1.600 3.180 1.645 ;
        RECT 0.550 1.460 3.180 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.890 1.415 3.180 1.460 ;
  END
END sky130_fd_sc_hd__dlxtn_2

#--------EOF---------

MACRO sky130_fd_sc_hd__dlxtn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.460 0.955 1.790 1.325 ;
    END
  END D
  PIN GATE_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.330 1.625 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 4.215 0.785 6.895 1.015 ;
        RECT 0.005 0.105 6.895 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER li1 ;
        RECT 5.240 1.495 5.525 2.455 ;
        RECT 5.355 1.325 5.525 1.495 ;
        RECT 6.115 1.325 6.385 2.455 ;
        RECT 5.355 0.995 6.815 1.325 ;
        RECT 5.355 0.745 5.525 0.995 ;
        RECT 5.240 0.415 5.525 0.745 ;
        RECT 6.115 0.385 6.385 0.995 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.175 0.635 0.780 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.455 1.665 1.785 2.415 ;
        RECT 1.955 1.835 2.270 2.635 ;
        RECT 2.900 2.255 3.650 2.425 ;
        RECT 1.455 1.495 2.140 1.665 ;
        RECT 1.970 1.095 2.140 1.495 ;
        RECT 2.470 1.355 2.755 2.005 ;
        RECT 2.925 1.415 3.265 1.995 ;
        RECT 1.970 0.785 2.340 1.095 ;
        RECT 2.925 1.035 3.095 1.415 ;
        RECT 3.480 1.325 3.650 2.255 ;
        RECT 3.820 2.135 4.120 2.635 ;
        RECT 4.385 1.865 4.605 2.435 ;
        RECT 3.840 1.535 4.605 1.865 ;
        RECT 4.435 1.325 4.605 1.535 ;
        RECT 4.785 1.495 5.070 2.635 ;
        RECT 5.695 1.495 5.945 2.635 ;
        RECT 6.555 1.495 6.815 2.635 ;
        RECT 3.480 1.165 4.200 1.325 ;
        RECT 1.535 0.765 2.340 0.785 ;
        RECT 1.535 0.615 2.140 0.765 ;
        RECT 2.715 0.705 3.095 1.035 ;
        RECT 3.330 0.995 4.200 1.165 ;
        RECT 4.435 0.995 5.185 1.325 ;
        RECT 1.535 0.345 1.705 0.615 ;
        RECT 3.330 0.535 3.500 0.995 ;
        RECT 4.435 0.745 4.605 0.995 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 2.840 0.365 3.500 0.535 ;
        RECT 3.740 0.085 4.070 0.530 ;
        RECT 4.385 0.415 4.605 0.745 ;
        RECT 4.785 0.085 5.070 0.715 ;
        RECT 5.695 0.085 5.945 0.825 ;
        RECT 6.555 0.085 6.815 0.715 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.470 1.785 2.640 1.955 ;
        RECT 2.930 1.445 3.100 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.410 1.940 2.700 1.985 ;
        RECT 1.010 1.800 2.700 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.410 1.755 2.700 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.870 1.600 3.160 1.645 ;
        RECT 0.550 1.460 3.160 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.870 1.415 3.160 1.460 ;
  END
END sky130_fd_sc_hd__dlxtn_4

#--------EOF---------

MACRO sky130_fd_sc_hd__dlxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.460 0.955 1.790 1.325 ;
    END
  END D
  PIN GATE
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.985 0.330 1.625 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.725 2.705 0.785 ;
        RECT 4.125 0.725 5.515 1.015 ;
        RECT 0.005 0.105 5.515 0.725 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER li1 ;
        RECT 5.150 1.670 5.435 2.455 ;
        RECT 5.265 0.745 5.435 1.670 ;
        RECT 5.150 0.415 5.435 0.745 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.610 1.400 0.780 1.795 ;
        RECT 1.015 1.685 1.240 2.465 ;
        RECT 0.610 1.070 0.840 1.400 ;
        RECT 0.610 0.805 0.780 1.070 ;
        RECT 0.175 0.635 0.780 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 1.685 ;
        RECT 1.455 1.665 1.785 2.415 ;
        RECT 1.955 1.835 2.270 2.635 ;
        RECT 2.770 2.255 3.605 2.425 ;
        RECT 1.455 1.495 2.140 1.665 ;
        RECT 1.970 1.095 2.140 1.495 ;
        RECT 2.470 1.355 2.755 1.685 ;
        RECT 2.925 1.575 3.265 1.995 ;
        RECT 1.970 0.785 2.340 1.095 ;
        RECT 2.925 1.035 3.095 1.575 ;
        RECT 3.435 1.325 3.605 2.255 ;
        RECT 3.775 2.135 3.945 2.635 ;
        RECT 4.295 1.865 4.515 2.435 ;
        RECT 3.840 1.535 4.515 1.865 ;
        RECT 4.695 1.570 4.900 2.635 ;
        RECT 4.345 1.325 4.515 1.535 ;
        RECT 3.435 1.165 4.175 1.325 ;
        RECT 1.535 0.765 2.340 0.785 ;
        RECT 1.535 0.615 2.140 0.765 ;
        RECT 2.715 0.705 3.095 1.035 ;
        RECT 3.330 0.995 4.175 1.165 ;
        RECT 4.345 0.995 5.095 1.325 ;
        RECT 1.535 0.345 1.705 0.615 ;
        RECT 3.330 0.535 3.500 0.995 ;
        RECT 4.345 0.745 4.515 0.995 ;
        RECT 1.875 0.085 2.205 0.445 ;
        RECT 2.840 0.365 3.500 0.535 ;
        RECT 3.685 0.085 4.015 0.530 ;
        RECT 4.295 0.415 4.515 0.745 ;
        RECT 4.695 0.085 4.900 0.715 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.610 1.445 0.780 1.615 ;
        RECT 1.070 1.785 1.240 1.955 ;
        RECT 2.930 1.785 3.100 1.955 ;
        RECT 2.470 1.445 2.640 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
      LAYER met1 ;
        RECT 1.010 1.940 1.300 1.985 ;
        RECT 2.870 1.940 3.160 1.985 ;
        RECT 1.010 1.800 3.160 1.940 ;
        RECT 1.010 1.755 1.300 1.800 ;
        RECT 2.870 1.755 3.160 1.800 ;
        RECT 0.550 1.600 0.840 1.645 ;
        RECT 2.410 1.600 2.700 1.645 ;
        RECT 0.550 1.460 2.700 1.600 ;
        RECT 0.550 1.415 0.840 1.460 ;
        RECT 2.410 1.415 2.700 1.460 ;
  END
END sky130_fd_sc_hd__dlxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dlygate4sd1_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlygate4sd1_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.555 1.615 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.365 0.785 2.780 1.015 ;
        RECT 0.005 0.105 2.780 0.785 ;
        RECT 0.140 -0.085 0.310 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 2.440 1.495 2.700 2.465 ;
        RECT 2.530 0.825 2.700 1.495 ;
        RECT 2.410 0.255 2.700 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 2.005 0.380 2.465 ;
        RECT 0.550 2.175 0.765 2.635 ;
        RECT 0.935 2.175 1.320 2.465 ;
        RECT 0.085 1.785 0.895 2.005 ;
        RECT 0.725 1.325 0.895 1.785 ;
        RECT 0.725 0.995 0.980 1.325 ;
        RECT 1.150 1.275 1.320 2.175 ;
        RECT 1.515 1.745 1.740 2.430 ;
        RECT 1.910 1.915 2.270 2.635 ;
        RECT 1.515 1.575 2.240 1.745 ;
        RECT 2.070 1.325 2.240 1.575 ;
        RECT 1.150 1.075 1.900 1.275 ;
        RECT 0.725 0.885 0.895 0.995 ;
        RECT 0.095 0.715 0.895 0.885 ;
        RECT 0.095 0.255 0.380 0.715 ;
        RECT 1.150 0.545 1.320 1.075 ;
        RECT 2.070 0.995 2.360 1.325 ;
        RECT 2.070 0.905 2.240 0.995 ;
        RECT 0.550 0.085 0.765 0.545 ;
        RECT 0.935 0.255 1.320 0.545 ;
        RECT 1.515 0.735 2.240 0.905 ;
        RECT 1.515 0.255 1.740 0.735 ;
        RECT 1.910 0.085 2.240 0.565 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__dlygate4sd1_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dlygate4sd2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlygate4sd2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.625 1.615 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.020 0.785 2.940 1.015 ;
        RECT 0.115 0.105 2.940 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 2.570 1.495 3.135 2.465 ;
        RECT 2.675 0.825 3.135 1.495 ;
        RECT 2.570 0.255 3.135 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 2.005 0.485 2.465 ;
        RECT 0.655 2.175 0.925 2.635 ;
        RECT 1.155 2.135 1.425 2.465 ;
        RECT 0.085 1.785 1.030 2.005 ;
        RECT 0.795 1.325 1.030 1.785 ;
        RECT 1.255 1.615 1.425 2.135 ;
        RECT 1.615 2.005 1.875 2.465 ;
        RECT 2.075 2.175 2.400 2.635 ;
        RECT 1.615 1.785 2.400 2.005 ;
        RECT 0.795 0.995 1.085 1.325 ;
        RECT 1.255 1.055 2.030 1.615 ;
        RECT 2.200 1.325 2.400 1.785 ;
        RECT 0.795 0.885 1.030 0.995 ;
        RECT 0.085 0.715 1.030 0.885 ;
        RECT 0.085 0.255 0.485 0.715 ;
        RECT 1.255 0.585 1.425 1.055 ;
        RECT 2.200 0.995 2.505 1.325 ;
        RECT 2.200 0.885 2.400 0.995 ;
        RECT 0.655 0.085 0.925 0.545 ;
        RECT 1.155 0.255 1.425 0.585 ;
        RECT 1.615 0.715 2.400 0.885 ;
        RECT 1.615 0.255 1.875 0.715 ;
        RECT 2.075 0.085 2.400 0.545 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__dlygate4sd2_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dlygate4sd3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlygate4sd3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 0.775 1.615 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.660 0.785 3.580 1.015 ;
        RECT 0.115 0.105 3.580 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 3.210 1.495 3.595 2.465 ;
        RECT 3.315 0.825 3.595 1.495 ;
        RECT 3.210 0.255 3.595 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.200 2.005 0.485 2.465 ;
        RECT 0.655 2.175 0.925 2.635 ;
        RECT 0.200 1.785 1.155 2.005 ;
        RECT 0.945 0.885 1.155 1.785 ;
        RECT 0.200 0.715 1.155 0.885 ;
        RECT 1.325 1.615 1.725 2.465 ;
        RECT 1.915 2.005 2.195 2.465 ;
        RECT 2.715 2.175 3.040 2.635 ;
        RECT 1.915 1.785 3.040 2.005 ;
        RECT 1.325 1.055 2.420 1.615 ;
        RECT 2.590 1.325 3.040 1.785 ;
        RECT 0.200 0.255 0.485 0.715 ;
        RECT 0.655 0.085 0.925 0.545 ;
        RECT 1.325 0.255 1.725 1.055 ;
        RECT 2.590 0.995 3.145 1.325 ;
        RECT 2.590 0.885 3.040 0.995 ;
        RECT 1.915 0.715 3.040 0.885 ;
        RECT 1.915 0.255 2.195 0.715 ;
        RECT 2.715 0.085 3.040 0.545 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__dlygate4sd3_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dlymetal6s2s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlymetal6s2s_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.570 1.700 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.665 0.785 4.595 1.015 ;
        RECT 0.180 0.105 4.595 0.785 ;
        RECT 0.180 0.085 0.290 0.105 ;
        RECT 0.120 -0.085 0.290 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 1.245 1.675 1.670 2.465 ;
        RECT 1.245 1.495 2.150 1.675 ;
        RECT 1.320 0.995 2.150 1.495 ;
        RECT 1.320 0.825 1.670 0.995 ;
        RECT 1.245 0.255 1.670 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.085 2.040 0.520 2.465 ;
        RECT 0.690 2.210 1.075 2.635 ;
        RECT 1.840 2.040 2.115 2.465 ;
        RECT 2.285 2.210 2.670 2.635 ;
        RECT 0.085 1.870 1.075 2.040 ;
        RECT 0.740 1.325 1.075 1.870 ;
        RECT 1.840 1.845 2.670 2.040 ;
        RECT 2.320 1.325 2.670 1.845 ;
        RECT 2.840 1.675 3.085 2.465 ;
        RECT 3.275 2.040 3.530 2.465 ;
        RECT 3.700 2.210 4.085 2.635 ;
        RECT 3.275 1.845 4.085 2.040 ;
        RECT 2.840 1.495 3.565 1.675 ;
        RECT 0.740 0.995 1.150 1.325 ;
        RECT 2.320 0.995 2.745 1.325 ;
        RECT 2.915 0.995 3.565 1.495 ;
        RECT 3.735 1.325 4.085 1.845 ;
        RECT 4.255 1.495 4.515 2.465 ;
        RECT 3.735 0.995 4.160 1.325 ;
        RECT 0.740 0.825 1.075 0.995 ;
        RECT 2.320 0.825 2.670 0.995 ;
        RECT 2.915 0.825 3.085 0.995 ;
        RECT 3.735 0.825 4.085 0.995 ;
        RECT 4.330 0.825 4.515 1.495 ;
        RECT 0.085 0.655 1.075 0.825 ;
        RECT 1.860 0.655 2.670 0.825 ;
        RECT 0.085 0.255 0.520 0.655 ;
        RECT 0.690 0.085 1.075 0.485 ;
        RECT 1.860 0.255 2.115 0.655 ;
        RECT 2.285 0.085 2.670 0.485 ;
        RECT 2.840 0.255 3.085 0.825 ;
        RECT 3.275 0.655 4.085 0.825 ;
        RECT 3.275 0.255 3.530 0.655 ;
        RECT 3.700 0.085 4.085 0.485 ;
        RECT 4.255 0.255 4.515 0.825 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__dlymetal6s2s_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dlymetal6s4s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlymetal6s4s_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.570 1.700 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.665 0.785 4.595 1.015 ;
        RECT 0.180 0.105 4.595 0.785 ;
        RECT 0.180 0.085 0.290 0.105 ;
        RECT 0.120 -0.085 0.290 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 2.660 1.675 3.105 2.465 ;
        RECT 2.660 1.495 3.565 1.675 ;
        RECT 2.735 0.995 3.565 1.495 ;
        RECT 2.735 0.825 3.105 0.995 ;
        RECT 2.660 0.255 3.105 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.085 2.040 0.520 2.465 ;
        RECT 0.690 2.210 1.075 2.635 ;
        RECT 0.085 1.870 1.075 2.040 ;
        RECT 0.740 1.325 1.075 1.870 ;
        RECT 1.245 1.675 1.515 2.465 ;
        RECT 1.685 2.040 1.935 2.465 ;
        RECT 2.105 2.210 2.490 2.635 ;
        RECT 3.275 2.040 3.530 2.465 ;
        RECT 3.700 2.210 4.085 2.635 ;
        RECT 1.685 1.845 2.490 2.040 ;
        RECT 3.275 1.845 4.085 2.040 ;
        RECT 1.245 1.495 1.970 1.675 ;
        RECT 0.740 0.995 1.150 1.325 ;
        RECT 1.320 0.995 1.970 1.495 ;
        RECT 2.140 1.325 2.490 1.845 ;
        RECT 3.735 1.325 4.085 1.845 ;
        RECT 4.255 1.495 4.515 2.465 ;
        RECT 2.140 0.995 2.565 1.325 ;
        RECT 3.735 0.995 4.160 1.325 ;
        RECT 0.740 0.825 1.075 0.995 ;
        RECT 1.320 0.825 1.515 0.995 ;
        RECT 2.140 0.825 2.490 0.995 ;
        RECT 3.735 0.825 4.085 0.995 ;
        RECT 4.330 0.825 4.515 1.495 ;
        RECT 0.085 0.655 1.075 0.825 ;
        RECT 0.085 0.255 0.520 0.655 ;
        RECT 0.690 0.085 1.075 0.485 ;
        RECT 1.245 0.255 1.515 0.825 ;
        RECT 1.685 0.655 2.490 0.825 ;
        RECT 3.275 0.655 4.085 0.825 ;
        RECT 1.685 0.255 1.935 0.655 ;
        RECT 2.105 0.085 2.490 0.485 ;
        RECT 3.275 0.255 3.530 0.655 ;
        RECT 3.700 0.085 4.085 0.485 ;
        RECT 4.255 0.255 4.515 0.825 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__dlymetal6s4s_1

#--------EOF---------

MACRO sky130_fd_sc_hd__dlymetal6s6s_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__dlymetal6s6s_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.575 1.700 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.670 0.785 4.420 1.015 ;
        RECT 0.185 0.105 4.420 0.785 ;
        RECT 0.185 0.085 0.295 0.105 ;
        RECT 0.125 -0.085 0.295 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 4.080 1.495 4.515 2.465 ;
        RECT 4.155 0.825 4.515 1.495 ;
        RECT 4.080 0.255 4.515 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.085 2.040 0.525 2.465 ;
        RECT 0.695 2.210 1.080 2.635 ;
        RECT 0.085 1.870 1.080 2.040 ;
        RECT 0.745 1.325 1.080 1.870 ;
        RECT 1.250 1.675 1.520 2.465 ;
        RECT 1.690 2.040 1.940 2.465 ;
        RECT 2.110 2.210 2.495 2.635 ;
        RECT 1.690 1.845 2.495 2.040 ;
        RECT 1.250 1.495 1.975 1.675 ;
        RECT 0.745 0.995 1.155 1.325 ;
        RECT 1.325 0.995 1.975 1.495 ;
        RECT 2.145 1.325 2.495 1.845 ;
        RECT 2.665 1.675 2.915 2.465 ;
        RECT 3.085 2.040 3.355 2.465 ;
        RECT 3.525 2.210 3.910 2.635 ;
        RECT 3.085 1.845 3.910 2.040 ;
        RECT 2.665 1.495 3.390 1.675 ;
        RECT 2.145 0.995 2.570 1.325 ;
        RECT 2.740 0.995 3.390 1.495 ;
        RECT 3.560 1.325 3.910 1.845 ;
        RECT 3.560 0.995 3.985 1.325 ;
        RECT 0.745 0.825 1.080 0.995 ;
        RECT 1.325 0.825 1.520 0.995 ;
        RECT 2.145 0.825 2.495 0.995 ;
        RECT 2.740 0.825 2.915 0.995 ;
        RECT 3.560 0.825 3.910 0.995 ;
        RECT 0.085 0.655 1.080 0.825 ;
        RECT 0.085 0.255 0.525 0.655 ;
        RECT 0.695 0.085 1.080 0.485 ;
        RECT 1.250 0.255 1.520 0.825 ;
        RECT 1.690 0.655 2.495 0.825 ;
        RECT 1.690 0.255 1.940 0.655 ;
        RECT 2.110 0.085 2.495 0.485 ;
        RECT 2.665 0.255 2.915 0.825 ;
        RECT 3.085 0.655 3.910 0.825 ;
        RECT 3.085 0.255 3.355 0.655 ;
        RECT 3.525 0.085 3.910 0.485 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__dlymetal6s6s_1

#--------EOF---------

MACRO sky130_fd_sc_hd__ebufn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.355 1.615 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.309000 ;
    PORT
      LAYER li1 ;
        RECT 0.910 1.075 1.240 1.630 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.490 0.785 3.585 1.015 ;
        RECT 0.005 0.335 3.585 0.785 ;
        RECT 0.005 0.105 0.955 0.335 ;
        RECT 2.025 0.105 3.585 0.335 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.601000 ;
    PORT
      LAYER li1 ;
        RECT 1.975 1.495 3.595 2.465 ;
        RECT 3.255 0.825 3.595 1.495 ;
        RECT 3.125 0.255 3.595 0.825 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 2.005 0.345 2.465 ;
        RECT 0.515 2.175 0.845 2.635 ;
        RECT 1.015 2.005 1.270 2.460 ;
        RECT 1.440 2.175 1.805 2.635 ;
        RECT 0.085 1.785 0.740 2.005 ;
        RECT 1.015 1.800 1.805 2.005 ;
        RECT 0.525 0.825 0.740 1.785 ;
        RECT 1.410 1.325 1.805 1.800 ;
        RECT 1.410 1.075 2.535 1.325 ;
        RECT 1.410 0.885 1.685 1.075 ;
        RECT 2.705 0.995 3.085 1.325 ;
        RECT 2.705 0.905 2.955 0.995 ;
        RECT 0.085 0.615 1.185 0.825 ;
        RECT 1.355 0.635 1.685 0.885 ;
        RECT 1.855 0.735 2.955 0.905 ;
        RECT 0.085 0.280 0.345 0.615 ;
        RECT 1.015 0.465 1.185 0.615 ;
        RECT 1.855 0.465 2.025 0.735 ;
        RECT 0.515 0.085 0.845 0.445 ;
        RECT 1.015 0.255 2.025 0.465 ;
        RECT 2.195 0.085 2.955 0.565 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__ebufn_1

#--------EOF---------

MACRO sky130_fd_sc_hd__ebufn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.490 0.765 0.780 1.675 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.441000 ;
    PORT
      LAYER li1 ;
        RECT 0.950 0.765 1.280 1.275 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.830 0.785 4.135 1.015 ;
        RECT 0.005 0.105 4.135 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 3.295 1.765 3.625 2.125 ;
        RECT 1.905 1.625 3.625 1.765 ;
        RECT 1.905 1.445 4.055 1.625 ;
        RECT 3.825 0.855 4.055 1.445 ;
        RECT 3.295 0.635 4.055 0.855 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 1.845 0.345 2.465 ;
        RECT 0.515 1.845 0.950 2.635 ;
        RECT 0.085 0.615 0.320 1.845 ;
        RECT 1.120 1.765 1.410 2.465 ;
        RECT 1.600 2.105 1.810 2.465 ;
        RECT 1.980 2.275 2.310 2.635 ;
        RECT 2.480 2.295 4.055 2.465 ;
        RECT 2.480 2.105 3.125 2.295 ;
        RECT 1.600 1.935 3.125 2.105 ;
        RECT 3.795 1.795 4.055 2.295 ;
        RECT 1.120 1.445 1.735 1.765 ;
        RECT 1.450 1.275 1.735 1.445 ;
        RECT 1.450 1.025 2.965 1.275 ;
        RECT 3.245 1.025 3.655 1.275 ;
        RECT 0.085 0.280 0.345 0.615 ;
        RECT 1.450 0.595 1.730 1.025 ;
        RECT 0.515 0.085 0.850 0.595 ;
        RECT 1.020 0.255 1.730 0.595 ;
        RECT 1.900 0.655 3.125 0.855 ;
        RECT 1.900 0.255 2.170 0.655 ;
        RECT 2.340 0.085 2.670 0.485 ;
        RECT 2.840 0.465 3.125 0.655 ;
        RECT 2.840 0.275 4.050 0.465 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.150 1.105 0.320 1.275 ;
        RECT 3.380 1.105 3.550 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
      LAYER met1 ;
        RECT 0.085 1.260 0.380 1.305 ;
        RECT 3.320 1.260 3.610 1.305 ;
        RECT 0.085 1.120 3.610 1.260 ;
        RECT 0.085 1.075 0.380 1.120 ;
        RECT 3.320 1.075 3.610 1.120 ;
  END
END sky130_fd_sc_hd__ebufn_2

#--------EOF---------

MACRO sky130_fd_sc_hd__ebufn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.490 0.765 0.780 1.675 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.811500 ;
    PORT
      LAYER li1 ;
        RECT 0.950 0.765 1.280 1.425 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.845 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 1.895 1.445 5.895 1.725 ;
        RECT 5.675 0.855 5.895 1.445 ;
        RECT 4.145 0.615 5.895 0.855 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.085 1.765 0.345 2.465 ;
        RECT 0.515 1.845 0.930 2.635 ;
        RECT 1.100 1.765 1.355 2.465 ;
        RECT 1.565 2.105 1.810 2.465 ;
        RECT 1.980 2.275 2.310 2.635 ;
        RECT 2.480 2.105 2.650 2.465 ;
        RECT 2.820 2.275 3.150 2.635 ;
        RECT 3.320 2.105 5.895 2.465 ;
        RECT 1.565 1.935 5.895 2.105 ;
        RECT 1.895 1.895 5.895 1.935 ;
        RECT 0.085 0.665 0.320 1.765 ;
        RECT 1.100 1.595 1.725 1.765 ;
        RECT 1.450 1.275 1.725 1.595 ;
        RECT 1.450 1.025 3.810 1.275 ;
        RECT 3.980 1.025 5.505 1.275 ;
        RECT 0.085 0.280 0.345 0.665 ;
        RECT 1.450 0.595 1.725 1.025 ;
        RECT 0.515 0.085 0.930 0.595 ;
        RECT 1.100 0.255 1.725 0.595 ;
        RECT 1.895 0.655 3.975 0.855 ;
        RECT 1.895 0.255 2.175 0.655 ;
        RECT 2.345 0.085 2.675 0.485 ;
        RECT 2.845 0.275 3.015 0.655 ;
        RECT 3.185 0.085 3.515 0.485 ;
        RECT 3.685 0.445 3.975 0.655 ;
        RECT 3.685 0.255 5.735 0.445 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.150 1.105 0.320 1.275 ;
        RECT 4.310 1.105 4.480 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
      LAYER met1 ;
        RECT 0.085 1.260 0.380 1.305 ;
        RECT 4.250 1.260 4.540 1.305 ;
        RECT 0.085 1.120 4.540 1.260 ;
        RECT 0.085 1.075 0.380 1.120 ;
        RECT 4.250 1.075 4.540 1.120 ;
  END
END sky130_fd_sc_hd__ebufn_4

#--------EOF---------

MACRO sky130_fd_sc_hd__ebufn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ebufn_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.430 1.615 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.375500 ;
    PORT
      LAYER li1 ;
        RECT 0.970 1.325 1.305 1.695 ;
        RECT 0.970 0.995 1.430 1.325 ;
        RECT 0.970 0.620 1.305 0.995 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.655 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 1.995 1.445 9.575 1.725 ;
        RECT 9.325 0.855 9.575 1.445 ;
        RECT 6.275 0.615 9.575 0.855 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.085 1.785 0.445 2.635 ;
        RECT 0.615 1.615 0.800 2.465 ;
        RECT 0.970 1.865 1.305 2.635 ;
        RECT 0.600 0.995 0.800 1.615 ;
        RECT 1.475 1.495 1.825 2.465 ;
        RECT 1.995 2.065 2.245 2.465 ;
        RECT 2.415 2.235 2.745 2.635 ;
        RECT 2.915 2.065 3.085 2.465 ;
        RECT 3.255 2.235 3.585 2.635 ;
        RECT 3.755 2.065 3.925 2.465 ;
        RECT 4.095 2.235 4.425 2.635 ;
        RECT 4.595 2.065 4.765 2.465 ;
        RECT 4.935 2.235 5.265 2.635 ;
        RECT 5.435 2.065 9.575 2.465 ;
        RECT 1.995 1.895 9.575 2.065 ;
        RECT 0.085 0.085 0.445 0.825 ;
        RECT 0.615 0.280 0.800 0.995 ;
        RECT 1.600 1.275 1.825 1.495 ;
        RECT 1.600 1.025 5.925 1.275 ;
        RECT 6.175 1.025 9.155 1.275 ;
        RECT 1.600 0.825 1.985 1.025 ;
        RECT 0.970 0.085 1.305 0.445 ;
        RECT 1.475 0.255 1.985 0.825 ;
        RECT 2.155 0.655 6.105 0.855 ;
        RECT 2.155 0.255 2.485 0.655 ;
        RECT 2.655 0.085 2.985 0.485 ;
        RECT 3.155 0.275 3.325 0.655 ;
        RECT 3.495 0.085 3.825 0.485 ;
        RECT 3.995 0.255 4.165 0.655 ;
        RECT 4.335 0.085 4.665 0.485 ;
        RECT 4.835 0.275 5.005 0.655 ;
        RECT 5.175 0.085 5.505 0.485 ;
        RECT 5.675 0.445 6.105 0.655 ;
        RECT 5.675 0.255 9.575 0.445 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.605 1.105 0.775 1.275 ;
        RECT 6.580 1.105 6.750 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 0.545 1.260 0.835 1.305 ;
        RECT 6.520 1.260 6.810 1.305 ;
        RECT 0.545 1.120 6.810 1.260 ;
        RECT 0.545 1.075 0.835 1.120 ;
        RECT 6.520 1.075 6.810 1.120 ;
  END
END sky130_fd_sc_hd__ebufn_8

#--------EOF---------

MACRO sky130_fd_sc_hd__edfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__edfxbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.960 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.720 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 2.110 1.185 2.325 1.370 ;
        RECT 2.110 0.765 2.565 1.185 ;
    END
  END DE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.960 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.100 0.785 7.020 1.005 ;
        RECT 9.005 0.785 11.655 1.015 ;
        RECT 0.005 0.725 4.545 0.785 ;
        RECT 5.505 0.725 11.655 0.785 ;
        RECT 0.005 0.105 11.655 0.725 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.150 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.960 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER li1 ;
        RECT 11.225 0.255 11.555 2.420 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 9.400 1.410 9.730 2.465 ;
        RECT 9.400 1.065 9.845 1.410 ;
        RECT 9.515 0.255 9.845 1.065 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.960 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.845 1.965 ;
        RECT 0.615 0.805 0.845 1.795 ;
        RECT 0.175 0.635 0.845 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 2.465 ;
        RECT 1.355 1.890 1.785 2.465 ;
        RECT 2.235 1.890 2.565 2.635 ;
        RECT 1.355 0.515 1.525 1.890 ;
        RECT 2.755 1.720 3.085 2.425 ;
        RECT 3.265 1.825 3.460 2.635 ;
        RECT 4.125 2.020 4.455 2.465 ;
        RECT 4.915 2.175 5.955 2.375 ;
        RECT 4.125 1.820 4.515 2.020 ;
        RECT 2.495 1.355 3.085 1.720 ;
        RECT 2.780 1.175 3.085 1.355 ;
        RECT 3.805 1.320 4.175 1.650 ;
        RECT 2.780 0.845 3.635 1.175 ;
        RECT 1.355 0.255 1.785 0.515 ;
        RECT 2.235 0.085 2.565 0.515 ;
        RECT 2.780 0.255 3.005 0.845 ;
        RECT 3.805 0.685 3.975 1.320 ;
        RECT 4.345 1.150 4.515 1.820 ;
        RECT 4.145 0.980 4.515 1.150 ;
        RECT 4.795 1.125 4.980 1.720 ;
        RECT 5.150 1.655 5.615 2.005 ;
        RECT 3.185 0.085 3.515 0.610 ;
        RECT 4.145 0.255 4.415 0.980 ;
        RECT 5.150 0.955 5.320 1.655 ;
        RECT 5.785 1.575 5.955 2.175 ;
        RECT 6.125 1.835 6.360 2.635 ;
        RECT 5.785 1.485 6.360 1.575 ;
        RECT 4.815 0.735 5.320 0.955 ;
        RECT 5.510 1.315 6.360 1.485 ;
        RECT 5.510 0.565 5.680 1.315 ;
        RECT 6.190 1.245 6.360 1.315 ;
        RECT 6.530 1.375 6.860 2.465 ;
        RECT 7.070 2.105 7.360 2.635 ;
        RECT 7.925 2.165 8.890 2.355 ;
        RECT 5.870 1.065 6.070 1.095 ;
        RECT 6.530 1.065 7.445 1.375 ;
        RECT 7.790 1.245 7.980 1.965 ;
        RECT 5.870 1.045 7.445 1.065 ;
        RECT 5.870 0.765 6.935 1.045 ;
        RECT 8.150 1.035 8.470 1.995 ;
        RECT 5.005 0.255 5.680 0.565 ;
        RECT 5.945 0.085 6.340 0.560 ;
        RECT 6.530 0.255 6.935 0.765 ;
        RECT 8.005 0.705 8.470 1.035 ;
        RECT 7.165 0.085 7.440 0.615 ;
        RECT 8.640 0.535 8.890 2.165 ;
        RECT 9.060 1.495 9.230 2.635 ;
        RECT 9.900 1.575 10.130 2.010 ;
        RECT 10.300 1.220 10.640 2.465 ;
        RECT 10.810 1.465 11.055 2.635 ;
        RECT 8.025 0.330 8.890 0.535 ;
        RECT 9.095 0.085 9.345 0.900 ;
        RECT 10.015 0.890 10.640 1.220 ;
        RECT 10.300 0.255 10.640 0.890 ;
        RECT 10.810 0.085 11.055 0.900 ;
        RECT 0.000 -0.085 11.960 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 0.635 1.785 0.805 1.955 ;
        RECT 1.015 1.445 1.185 1.615 ;
        RECT 1.355 0.425 1.525 0.595 ;
        RECT 5.210 1.785 5.380 1.955 ;
        RECT 3.805 0.765 3.975 0.935 ;
        RECT 4.800 1.445 4.970 1.615 ;
        RECT 4.185 0.425 4.355 0.595 ;
        RECT 7.800 1.785 7.970 1.955 ;
        RECT 8.220 1.445 8.390 1.615 ;
        RECT 8.680 1.785 8.850 1.955 ;
        RECT 9.930 1.785 10.100 1.955 ;
        RECT 10.390 0.765 10.560 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
      LAYER met1 ;
        RECT 0.575 1.940 0.865 1.985 ;
        RECT 5.150 1.940 5.440 1.985 ;
        RECT 7.740 1.940 8.030 1.985 ;
        RECT 0.575 1.800 8.030 1.940 ;
        RECT 0.575 1.755 0.865 1.800 ;
        RECT 5.150 1.755 5.440 1.800 ;
        RECT 7.740 1.755 8.030 1.800 ;
        RECT 8.620 1.940 8.910 1.985 ;
        RECT 9.870 1.940 10.160 1.985 ;
        RECT 8.620 1.800 10.160 1.940 ;
        RECT 8.620 1.755 8.910 1.800 ;
        RECT 9.870 1.755 10.160 1.800 ;
        RECT 0.955 1.600 1.245 1.645 ;
        RECT 4.740 1.600 5.030 1.645 ;
        RECT 8.160 1.600 8.450 1.645 ;
        RECT 0.955 1.460 8.450 1.600 ;
        RECT 0.955 1.415 1.245 1.460 ;
        RECT 4.740 1.415 5.030 1.460 ;
        RECT 8.160 1.415 8.450 1.460 ;
        RECT 3.745 0.920 4.035 0.965 ;
        RECT 10.330 0.920 10.620 0.965 ;
        RECT 3.745 0.780 10.620 0.920 ;
        RECT 3.745 0.735 4.035 0.780 ;
        RECT 10.330 0.735 10.620 0.780 ;
        RECT 1.295 0.580 1.585 0.625 ;
        RECT 4.125 0.580 4.415 0.625 ;
        RECT 1.295 0.395 4.415 0.580 ;
  END
END sky130_fd_sc_hd__edfxbp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__edfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__edfxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.720 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 2.110 1.185 2.325 1.370 ;
        RECT 2.110 0.765 2.565 1.185 ;
    END
  END DE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.100 0.785 7.020 1.005 ;
        RECT 9.945 0.785 10.895 1.015 ;
        RECT 0.005 0.725 4.545 0.785 ;
        RECT 5.505 0.725 10.895 0.785 ;
        RECT 0.005 0.105 10.895 0.725 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER li1 ;
        RECT 10.465 0.305 10.795 2.420 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.845 1.965 ;
        RECT 0.615 0.805 0.845 1.795 ;
        RECT 0.175 0.635 0.845 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 2.465 ;
        RECT 1.355 1.890 1.785 2.465 ;
        RECT 2.235 1.890 2.565 2.635 ;
        RECT 1.355 0.515 1.525 1.890 ;
        RECT 2.755 1.720 3.085 2.425 ;
        RECT 3.265 1.825 3.460 2.635 ;
        RECT 4.125 2.020 4.455 2.465 ;
        RECT 4.915 2.175 5.955 2.375 ;
        RECT 4.125 1.820 4.515 2.020 ;
        RECT 2.495 1.355 3.085 1.720 ;
        RECT 2.780 1.175 3.085 1.355 ;
        RECT 3.805 1.320 4.175 1.650 ;
        RECT 2.780 0.845 3.635 1.175 ;
        RECT 1.355 0.255 1.785 0.515 ;
        RECT 2.235 0.085 2.565 0.515 ;
        RECT 2.780 0.255 3.005 0.845 ;
        RECT 3.805 0.685 3.975 1.320 ;
        RECT 4.345 1.150 4.515 1.820 ;
        RECT 4.145 0.980 4.515 1.150 ;
        RECT 4.795 1.125 4.980 1.720 ;
        RECT 5.150 1.655 5.615 2.005 ;
        RECT 3.185 0.085 3.515 0.610 ;
        RECT 4.145 0.255 4.415 0.980 ;
        RECT 5.150 0.955 5.320 1.655 ;
        RECT 5.785 1.575 5.955 2.175 ;
        RECT 6.125 1.835 6.360 2.635 ;
        RECT 5.785 1.485 6.360 1.575 ;
        RECT 4.815 0.735 5.320 0.955 ;
        RECT 5.510 1.315 6.360 1.485 ;
        RECT 5.510 0.565 5.680 1.315 ;
        RECT 6.190 1.245 6.360 1.315 ;
        RECT 6.530 1.375 6.860 2.465 ;
        RECT 7.070 2.105 7.360 2.635 ;
        RECT 7.925 2.165 8.810 2.355 ;
        RECT 5.870 1.065 6.070 1.095 ;
        RECT 6.530 1.065 7.445 1.375 ;
        RECT 7.790 1.245 7.980 1.965 ;
        RECT 5.870 1.045 7.445 1.065 ;
        RECT 5.870 0.765 6.935 1.045 ;
        RECT 8.150 1.035 8.470 1.995 ;
        RECT 5.005 0.255 5.680 0.565 ;
        RECT 5.945 0.085 6.340 0.560 ;
        RECT 6.530 0.255 6.935 0.765 ;
        RECT 8.005 0.705 8.470 1.035 ;
        RECT 8.640 1.325 8.810 2.165 ;
        RECT 8.980 2.135 9.240 2.635 ;
        RECT 9.540 1.905 9.880 2.465 ;
        RECT 8.980 1.530 9.880 1.905 ;
        RECT 8.640 0.995 9.510 1.325 ;
        RECT 7.165 0.085 7.440 0.615 ;
        RECT 8.640 0.535 8.810 0.995 ;
        RECT 9.690 0.825 9.880 1.530 ;
        RECT 10.050 1.465 10.295 2.635 ;
        RECT 8.025 0.330 8.810 0.535 ;
        RECT 9.050 0.085 9.365 0.615 ;
        RECT 9.550 0.300 9.880 0.825 ;
        RECT 10.050 0.085 10.295 0.900 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 0.635 1.785 0.805 1.955 ;
        RECT 1.015 1.445 1.185 1.615 ;
        RECT 1.355 0.425 1.525 0.595 ;
        RECT 5.210 1.785 5.380 1.955 ;
        RECT 3.805 0.765 3.975 0.935 ;
        RECT 4.800 1.445 4.970 1.615 ;
        RECT 4.185 0.425 4.355 0.595 ;
        RECT 7.800 1.785 7.970 1.955 ;
        RECT 8.220 1.445 8.390 1.615 ;
        RECT 9.700 0.765 9.870 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
      LAYER met1 ;
        RECT 0.575 1.940 0.865 1.985 ;
        RECT 5.150 1.940 5.440 1.985 ;
        RECT 7.740 1.940 8.030 1.985 ;
        RECT 0.575 1.800 8.030 1.940 ;
        RECT 0.575 1.755 0.865 1.800 ;
        RECT 5.150 1.755 5.440 1.800 ;
        RECT 7.740 1.755 8.030 1.800 ;
        RECT 0.955 1.600 1.245 1.645 ;
        RECT 4.740 1.600 5.030 1.645 ;
        RECT 8.160 1.600 8.450 1.645 ;
        RECT 0.955 1.460 8.450 1.600 ;
        RECT 0.955 1.415 1.245 1.460 ;
        RECT 4.740 1.415 5.030 1.460 ;
        RECT 8.160 1.415 8.450 1.460 ;
        RECT 3.745 0.920 4.035 0.965 ;
        RECT 9.640 0.920 9.930 0.965 ;
        RECT 3.745 0.780 9.930 0.920 ;
        RECT 3.745 0.735 4.035 0.780 ;
        RECT 9.640 0.735 9.930 0.780 ;
        RECT 1.295 0.580 1.585 0.625 ;
        RECT 4.125 0.580 4.415 0.625 ;
        RECT 1.295 0.395 4.415 0.580 ;
  END
END sky130_fd_sc_hd__edfxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__einvn_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.500 0.765 1.755 1.955 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.222000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.650 1.725 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.020 0.105 1.825 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.275600 ;
    PORT
      LAYER li1 ;
        RECT 1.160 2.125 1.755 2.465 ;
        RECT 1.160 0.595 1.330 2.125 ;
        RECT 1.160 0.255 1.755 0.595 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.085 2.065 0.400 2.465 ;
        RECT 0.570 2.235 0.990 2.635 ;
        RECT 0.085 1.895 0.990 2.065 ;
        RECT 0.820 0.825 0.990 1.895 ;
        RECT 0.085 0.655 0.990 0.825 ;
        RECT 0.085 0.255 0.360 0.655 ;
        RECT 0.530 0.085 0.990 0.485 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__einvn_0

#--------EOF---------

MACRO sky130_fd_sc_hd__einvn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.970 0.765 2.215 1.615 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.309000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.510 1.725 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.490 0.785 2.295 1.015 ;
        RECT 0.005 0.105 2.295 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 1.040 1.785 2.215 2.465 ;
        RECT 1.620 0.595 1.800 1.785 ;
        RECT 1.620 0.255 2.215 0.595 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.085 2.065 0.370 2.465 ;
        RECT 0.540 2.235 0.870 2.635 ;
        RECT 0.085 1.895 0.870 2.065 ;
        RECT 0.685 1.615 0.870 1.895 ;
        RECT 0.685 0.785 1.450 1.615 ;
        RECT 0.085 0.615 1.450 0.785 ;
        RECT 0.085 0.255 0.370 0.615 ;
        RECT 0.540 0.085 1.440 0.445 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__einvn_1

#--------EOF---------

MACRO sky130_fd_sc_hd__einvn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.785 1.075 3.135 1.275 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.441000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.325 1.385 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.940 0.785 3.205 1.015 ;
        RECT 0.005 0.105 3.205 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.694800 ;
    PORT
      LAYER li1 ;
        RECT 2.785 1.695 3.135 2.465 ;
        RECT 1.945 1.445 3.135 1.695 ;
        RECT 2.365 0.845 2.615 1.445 ;
        RECT 2.365 0.595 2.695 0.845 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.725 0.345 2.465 ;
        RECT 0.515 1.895 0.895 2.635 ;
        RECT 1.070 2.085 1.240 2.465 ;
        RECT 1.410 2.255 2.275 2.635 ;
        RECT 2.445 2.085 2.615 2.465 ;
        RECT 1.070 1.865 2.615 2.085 ;
        RECT 0.085 1.555 0.895 1.725 ;
        RECT 0.495 1.275 0.895 1.555 ;
        RECT 1.070 1.445 1.775 1.865 ;
        RECT 0.495 0.995 2.035 1.275 ;
        RECT 0.495 0.825 0.840 0.995 ;
        RECT 0.085 0.655 0.840 0.825 ;
        RECT 1.015 0.655 2.195 0.825 ;
        RECT 0.085 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.015 0.255 1.280 0.655 ;
        RECT 1.450 0.085 1.780 0.485 ;
        RECT 1.950 0.425 2.195 0.655 ;
        RECT 2.865 0.425 3.135 0.775 ;
        RECT 1.950 0.255 3.135 0.425 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__einvn_2

#--------EOF---------

MACRO sky130_fd_sc_hd__einvn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 4.530 0.620 4.975 1.325 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.811500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.345 1.325 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.890 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 3.190 1.480 3.520 2.075 ;
        RECT 4.030 1.480 4.360 2.075 ;
        RECT 3.190 0.620 4.360 1.480 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.085 1.665 0.345 2.465 ;
        RECT 0.515 1.835 0.845 2.635 ;
        RECT 1.015 1.665 1.240 2.465 ;
        RECT 1.410 1.835 1.740 2.635 ;
        RECT 1.910 1.665 2.080 2.465 ;
        RECT 2.250 1.835 2.640 2.635 ;
        RECT 2.810 2.295 4.975 2.465 ;
        RECT 2.810 1.665 3.020 2.295 ;
        RECT 0.085 1.495 0.845 1.665 ;
        RECT 1.015 1.495 3.020 1.665 ;
        RECT 3.690 1.650 3.860 2.295 ;
        RECT 4.530 1.650 4.975 2.295 ;
        RECT 0.515 1.325 0.845 1.495 ;
        RECT 0.515 0.995 3.020 1.325 ;
        RECT 0.515 0.825 0.845 0.995 ;
        RECT 0.085 0.655 0.845 0.825 ;
        RECT 1.015 0.655 2.995 0.825 ;
        RECT 0.085 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.015 0.255 1.285 0.655 ;
        RECT 1.455 0.085 1.785 0.485 ;
        RECT 1.955 0.255 2.125 0.655 ;
        RECT 2.295 0.085 2.625 0.485 ;
        RECT 2.825 0.450 2.995 0.655 ;
        RECT 2.825 0.255 4.975 0.450 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
END sky130_fd_sc_hd__einvn_4

#--------EOF---------

MACRO sky130_fd_sc_hd__einvn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvn_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 4.645 0.995 7.800 1.285 ;
    END
  END A
  PIN TE_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.375500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.995 0.345 1.325 ;
    END
  END TE_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.250 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 4.870 1.625 5.200 2.125 ;
        RECT 5.710 1.625 6.040 2.125 ;
        RECT 6.550 1.625 6.880 2.125 ;
        RECT 7.390 1.625 7.720 2.125 ;
        RECT 4.870 1.455 8.195 1.625 ;
        RECT 7.970 0.825 8.195 1.455 ;
        RECT 4.870 0.620 8.195 0.825 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.090 1.665 0.345 2.465 ;
        RECT 0.515 1.835 0.845 2.635 ;
        RECT 1.015 1.665 1.240 2.465 ;
        RECT 1.410 1.835 1.740 2.635 ;
        RECT 1.910 1.665 2.080 2.465 ;
        RECT 2.250 1.835 2.580 2.635 ;
        RECT 2.750 1.665 2.920 2.465 ;
        RECT 3.090 1.835 3.420 2.635 ;
        RECT 3.590 1.665 3.760 2.465 ;
        RECT 3.930 1.835 4.280 2.635 ;
        RECT 4.450 2.295 8.195 2.465 ;
        RECT 4.450 1.665 4.700 2.295 ;
        RECT 5.370 1.795 5.540 2.295 ;
        RECT 6.210 1.795 6.380 2.295 ;
        RECT 7.050 1.795 7.220 2.295 ;
        RECT 7.890 1.795 8.195 2.295 ;
        RECT 0.090 1.495 0.845 1.665 ;
        RECT 1.015 1.495 4.700 1.665 ;
        RECT 0.515 1.325 0.845 1.495 ;
        RECT 0.515 0.995 4.475 1.325 ;
        RECT 0.515 0.825 0.845 0.995 ;
        RECT 0.090 0.655 0.845 0.825 ;
        RECT 1.015 0.655 4.700 0.825 ;
        RECT 0.090 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.015 0.255 1.285 0.655 ;
        RECT 1.455 0.085 1.785 0.485 ;
        RECT 1.955 0.255 2.125 0.655 ;
        RECT 2.295 0.085 2.625 0.485 ;
        RECT 2.795 0.255 2.965 0.655 ;
        RECT 3.135 0.085 3.465 0.485 ;
        RECT 3.635 0.255 3.805 0.655 ;
        RECT 3.975 0.085 4.315 0.485 ;
        RECT 4.485 0.450 4.700 0.655 ;
        RECT 4.485 0.255 8.195 0.450 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
  END
END sky130_fd_sc_hd__einvn_8

#--------EOF---------

MACRO sky130_fd_sc_hd__einvp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.975 0.975 2.215 1.955 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.223500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.545 1.725 ;
    END
  END TE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.490 0.785 2.295 1.015 ;
        RECT 0.005 0.105 2.295 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 1.620 2.125 2.215 2.465 ;
        RECT 1.620 0.805 1.795 2.125 ;
        RECT 1.620 0.255 2.215 0.805 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.085 2.065 0.345 2.465 ;
        RECT 0.515 2.235 1.450 2.635 ;
        RECT 0.085 1.895 1.450 2.065 ;
        RECT 0.715 0.825 1.450 1.895 ;
        RECT 0.085 0.655 1.450 0.825 ;
        RECT 0.085 0.255 0.345 0.655 ;
        RECT 0.515 0.085 1.450 0.485 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__einvp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__einvp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.850 0.765 3.135 1.615 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.354000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.330 1.615 ;
    END
  END TE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.490 0.785 3.190 1.015 ;
        RECT 0.005 0.105 3.190 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 2.350 0.595 2.680 2.125 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.955 0.345 2.465 ;
        RECT 0.515 2.125 0.875 2.635 ;
        RECT 0.085 1.785 0.875 1.955 ;
        RECT 0.500 1.325 0.875 1.785 ;
        RECT 1.045 1.725 1.285 2.465 ;
        RECT 1.455 1.895 1.785 2.635 ;
        RECT 1.985 2.295 3.135 2.465 ;
        RECT 1.985 1.725 2.155 2.295 ;
        RECT 2.850 1.785 3.135 2.295 ;
        RECT 1.045 1.555 2.155 1.725 ;
        RECT 0.500 0.995 2.180 1.325 ;
        RECT 0.500 0.825 0.875 0.995 ;
        RECT 0.085 0.655 0.875 0.825 ;
        RECT 1.045 0.655 2.180 0.825 ;
        RECT 0.085 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.875 0.485 ;
        RECT 1.045 0.255 1.240 0.655 ;
        RECT 1.410 0.085 1.770 0.485 ;
        RECT 1.940 0.425 2.180 0.655 ;
        RECT 2.850 0.425 3.135 0.595 ;
        RECT 1.940 0.255 3.135 0.425 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__einvp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__einvp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.740 1.020 4.975 1.275 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.637500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.330 1.615 ;
    END
  END TE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.890 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 3.190 1.615 3.520 2.125 ;
        RECT 4.030 1.615 4.360 2.125 ;
        RECT 3.190 1.445 4.360 1.615 ;
        RECT 3.190 0.850 3.570 1.445 ;
        RECT 3.190 0.635 4.975 0.850 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.085 1.955 0.345 2.465 ;
        RECT 0.515 2.125 0.875 2.635 ;
        RECT 0.085 1.785 0.875 1.955 ;
        RECT 0.500 1.325 0.875 1.785 ;
        RECT 1.075 1.725 1.285 2.465 ;
        RECT 1.455 1.895 1.785 2.635 ;
        RECT 1.955 1.725 2.125 2.465 ;
        RECT 2.295 1.895 2.655 2.635 ;
        RECT 2.825 2.295 4.975 2.465 ;
        RECT 2.825 1.725 2.995 2.295 ;
        RECT 3.690 1.785 3.860 2.295 ;
        RECT 1.075 1.555 2.995 1.725 ;
        RECT 4.530 1.445 4.975 2.295 ;
        RECT 0.500 0.995 3.020 1.325 ;
        RECT 0.500 0.825 0.695 0.995 ;
        RECT 0.085 0.655 0.695 0.825 ;
        RECT 1.035 0.655 3.020 0.825 ;
        RECT 0.085 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.035 0.255 1.205 0.655 ;
        RECT 1.375 0.085 1.705 0.485 ;
        RECT 1.875 0.255 2.045 0.655 ;
        RECT 2.215 0.085 2.555 0.485 ;
        RECT 2.735 0.465 3.020 0.655 ;
        RECT 2.735 0.255 4.975 0.465 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
END sky130_fd_sc_hd__einvp_4

#--------EOF---------

MACRO sky130_fd_sc_hd__einvp_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__einvp_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 5.420 1.020 8.195 1.275 ;
    END
  END A
  PIN TE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.027500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.330 1.615 ;
    END
  END TE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.250 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 4.870 1.615 5.200 2.125 ;
        RECT 5.710 1.615 6.040 2.125 ;
        RECT 6.550 1.615 6.880 2.125 ;
        RECT 7.390 1.615 7.720 2.125 ;
        RECT 4.870 1.445 7.720 1.615 ;
        RECT 4.870 0.850 5.250 1.445 ;
        RECT 4.870 0.635 8.195 0.850 ;
    END
  END Z
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.085 1.955 0.345 2.465 ;
        RECT 0.515 2.125 0.875 2.635 ;
        RECT 0.085 1.785 0.875 1.955 ;
        RECT 0.500 1.325 0.875 1.785 ;
        RECT 1.075 1.725 1.285 2.465 ;
        RECT 1.455 1.895 1.785 2.635 ;
        RECT 1.955 1.725 2.125 2.465 ;
        RECT 2.295 1.895 2.625 2.635 ;
        RECT 2.795 1.725 2.965 2.465 ;
        RECT 3.135 1.895 3.465 2.635 ;
        RECT 3.635 1.725 3.805 2.465 ;
        RECT 3.975 1.895 4.305 2.635 ;
        RECT 4.475 2.295 8.195 2.465 ;
        RECT 4.475 1.725 4.700 2.295 ;
        RECT 5.370 1.785 5.540 2.295 ;
        RECT 6.210 1.785 6.380 2.295 ;
        RECT 7.050 1.785 7.220 2.295 ;
        RECT 1.075 1.555 4.700 1.725 ;
        RECT 7.890 1.445 8.195 2.295 ;
        RECT 0.500 0.995 4.700 1.325 ;
        RECT 0.500 0.825 0.695 0.995 ;
        RECT 0.085 0.655 0.695 0.825 ;
        RECT 1.035 0.655 4.700 0.825 ;
        RECT 0.085 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.035 0.255 1.205 0.655 ;
        RECT 1.375 0.085 1.705 0.485 ;
        RECT 1.875 0.255 2.045 0.655 ;
        RECT 2.215 0.085 2.545 0.485 ;
        RECT 2.715 0.255 2.885 0.655 ;
        RECT 3.055 0.085 3.385 0.485 ;
        RECT 3.555 0.255 3.725 0.655 ;
        RECT 3.895 0.085 4.235 0.485 ;
        RECT 4.405 0.465 4.700 0.655 ;
        RECT 4.405 0.255 8.195 0.465 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
  END
END sky130_fd_sc_hd__einvp_8

#--------EOF---------

MACRO sky130_fd_sc_hd__fa_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fa_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER met1 ;
        RECT 1.010 1.260 1.300 1.305 ;
        RECT 2.390 1.260 2.680 1.305 ;
        RECT 4.250 1.260 4.540 1.305 ;
        RECT 6.090 1.260 6.380 1.305 ;
        RECT 1.010 1.120 6.380 1.260 ;
        RECT 1.010 1.075 1.300 1.120 ;
        RECT 2.390 1.075 2.680 1.120 ;
        RECT 4.250 1.075 4.540 1.120 ;
        RECT 6.090 1.075 6.380 1.120 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER met1 ;
        RECT 1.470 1.600 1.760 1.645 ;
        RECT 3.330 1.600 3.620 1.645 ;
        RECT 5.630 1.600 5.920 1.645 ;
        RECT 1.470 1.460 5.920 1.600 ;
        RECT 1.470 1.415 1.760 1.460 ;
        RECT 3.330 1.415 3.620 1.460 ;
        RECT 5.630 1.415 5.920 1.460 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 1.870 1.595 2.960 1.765 ;
        RECT 5.155 1.685 5.405 1.955 ;
        RECT 1.870 1.275 2.040 1.595 ;
        RECT 1.670 1.105 2.040 1.275 ;
        RECT 2.790 1.250 2.960 1.595 ;
        RECT 3.785 1.515 5.405 1.685 ;
        RECT 3.785 1.250 3.955 1.515 ;
        RECT 2.790 0.965 3.955 1.250 ;
    END
  END CIN
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 0.935 1.015 ;
        RECT 6.250 0.785 7.180 1.015 ;
        RECT 0.005 0.105 7.180 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.485 0.345 2.465 ;
        RECT 0.085 0.830 0.260 1.485 ;
        RECT 0.085 0.255 0.345 0.830 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 6.840 1.485 7.240 2.465 ;
        RECT 6.910 0.810 7.240 1.485 ;
        RECT 6.840 0.255 7.240 0.810 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.515 2.150 0.765 2.635 ;
        RECT 0.935 2.065 1.710 2.465 ;
        RECT 1.960 2.105 2.130 2.465 ;
        RECT 2.300 2.275 2.630 2.635 ;
        RECT 2.800 2.105 3.035 2.465 ;
        RECT 3.240 2.255 3.570 2.635 ;
        RECT 0.935 1.945 1.105 2.065 ;
        RECT 0.515 1.625 1.105 1.945 ;
        RECT 1.960 1.935 3.035 2.105 ;
        RECT 3.740 2.105 3.910 2.465 ;
        RECT 4.080 2.275 4.410 2.635 ;
        RECT 4.580 2.105 4.750 2.465 ;
        RECT 5.085 2.125 6.170 2.465 ;
        RECT 6.340 2.275 6.670 2.635 ;
        RECT 3.740 1.935 4.750 2.105 ;
        RECT 6.000 2.105 6.170 2.125 ;
        RECT 6.000 1.935 6.665 2.105 ;
        RECT 0.515 1.325 0.685 1.625 ;
        RECT 1.300 1.445 1.700 1.880 ;
        RECT 3.200 1.435 3.560 1.765 ;
        RECT 5.635 1.445 6.055 1.765 ;
        RECT 0.430 0.995 0.685 1.325 ;
        RECT 0.910 1.275 1.080 1.325 ;
        RECT 0.910 0.995 1.240 1.275 ;
        RECT 2.230 1.030 2.620 1.360 ;
        RECT 6.495 1.325 6.665 1.935 ;
        RECT 0.515 0.805 0.685 0.995 ;
        RECT 4.250 0.955 4.625 1.275 ;
        RECT 4.795 0.955 5.460 1.125 ;
        RECT 5.885 1.035 6.325 1.275 ;
        RECT 1.470 0.805 1.710 0.935 ;
        RECT 0.515 0.635 1.710 0.805 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.110 0.255 1.710 0.635 ;
        RECT 1.960 0.615 2.970 0.785 ;
        RECT 1.960 0.255 2.130 0.615 ;
        RECT 2.300 0.085 2.630 0.445 ;
        RECT 2.800 0.255 2.970 0.615 ;
        RECT 3.740 0.615 4.750 0.785 ;
        RECT 4.965 0.765 5.460 0.955 ;
        RECT 6.495 0.995 6.740 1.325 ;
        RECT 6.495 0.785 6.665 0.995 ;
        RECT 3.240 0.085 3.570 0.490 ;
        RECT 3.740 0.255 3.910 0.615 ;
        RECT 4.080 0.085 4.410 0.445 ;
        RECT 4.580 0.255 4.750 0.615 ;
        RECT 5.925 0.615 6.665 0.785 ;
        RECT 5.085 0.505 5.255 0.595 ;
        RECT 5.925 0.505 6.095 0.615 ;
        RECT 5.085 0.255 6.095 0.505 ;
        RECT 6.265 0.085 6.595 0.445 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 1.530 1.445 1.700 1.615 ;
        RECT 3.390 1.445 3.560 1.615 ;
        RECT 5.690 1.445 5.860 1.615 ;
        RECT 1.070 1.105 1.240 1.275 ;
        RECT 2.450 1.105 2.620 1.275 ;
        RECT 4.310 1.105 4.480 1.275 ;
        RECT 6.150 1.105 6.320 1.275 ;
        RECT 1.530 0.765 1.700 0.935 ;
        RECT 5.230 0.765 5.400 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
      LAYER met1 ;
        RECT 1.470 0.920 1.760 0.965 ;
        RECT 5.170 0.920 5.460 0.965 ;
        RECT 1.470 0.780 5.460 0.920 ;
        RECT 1.470 0.735 1.760 0.780 ;
        RECT 5.170 0.735 5.460 0.780 ;
  END
END sky130_fd_sc_hd__fa_1

#--------EOF---------

MACRO sky130_fd_sc_hd__fa_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fa_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631500 ;
    PORT
      LAYER met1 ;
        RECT 1.465 1.260 1.755 1.305 ;
        RECT 2.845 1.260 3.135 1.305 ;
        RECT 4.705 1.260 4.995 1.305 ;
        RECT 6.085 1.260 6.375 1.305 ;
        RECT 1.465 1.120 6.375 1.260 ;
        RECT 1.465 1.075 1.755 1.120 ;
        RECT 2.845 1.075 3.135 1.120 ;
        RECT 4.705 1.075 4.995 1.120 ;
        RECT 6.085 1.075 6.375 1.120 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631500 ;
    PORT
      LAYER met1 ;
        RECT 1.925 1.600 2.215 1.645 ;
        RECT 3.785 1.600 4.075 1.645 ;
        RECT 6.545 1.600 6.835 1.645 ;
        RECT 1.925 1.460 6.835 1.600 ;
        RECT 1.925 1.415 2.215 1.460 ;
        RECT 3.785 1.415 4.075 1.460 ;
        RECT 6.545 1.415 6.835 1.460 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.475500 ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.570 3.415 1.740 ;
        RECT 5.670 1.685 5.920 1.955 ;
        RECT 2.325 1.275 2.495 1.570 ;
        RECT 2.125 1.105 2.495 1.275 ;
        RECT 3.245 1.250 3.415 1.570 ;
        RECT 4.295 1.515 5.920 1.685 ;
        RECT 4.295 1.435 4.655 1.515 ;
        RECT 4.295 1.250 4.465 1.435 ;
        RECT 5.670 1.355 5.920 1.515 ;
        RECT 3.245 0.965 4.465 1.250 ;
    END
  END CIN
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.785 1.360 1.015 ;
        RECT 6.765 0.785 8.235 1.015 ;
        RECT 0.010 0.105 8.235 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.600 1.950 0.810 2.465 ;
        RECT 0.565 1.780 0.810 1.950 ;
        RECT 0.565 1.585 0.735 1.780 ;
        RECT 0.085 1.415 0.735 1.585 ;
        RECT 0.085 0.905 0.370 1.415 ;
        RECT 0.085 0.735 0.690 0.905 ;
        RECT 0.520 0.485 0.690 0.735 ;
        RECT 0.520 0.315 0.850 0.485 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.523500 ;
    PORT
      LAYER li1 ;
        RECT 7.395 1.965 7.565 2.465 ;
        RECT 7.395 1.795 7.645 1.965 ;
        RECT 7.475 1.585 7.645 1.795 ;
        RECT 7.475 1.415 8.195 1.585 ;
        RECT 7.970 0.905 8.195 1.415 ;
        RECT 7.475 0.735 8.195 0.905 ;
        RECT 7.475 0.485 7.725 0.735 ;
        RECT 7.395 0.255 7.725 0.485 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.180 1.795 0.350 2.635 ;
        RECT 0.980 2.275 1.310 2.635 ;
        RECT 1.900 2.080 2.245 2.465 ;
        RECT 1.305 1.910 2.245 2.080 ;
        RECT 2.415 2.105 2.585 2.465 ;
        RECT 2.755 2.275 3.085 2.635 ;
        RECT 3.255 2.105 3.490 2.465 ;
        RECT 2.415 1.935 3.490 2.105 ;
        RECT 3.695 1.915 4.025 2.635 ;
        RECT 4.195 2.105 4.365 2.465 ;
        RECT 4.535 2.275 4.865 2.635 ;
        RECT 5.035 2.105 5.205 2.465 ;
        RECT 5.485 2.125 6.685 2.465 ;
        RECT 6.890 2.275 7.220 2.635 ;
        RECT 4.195 1.935 5.205 2.105 ;
        RECT 6.515 2.105 6.685 2.125 ;
        RECT 6.515 1.935 7.180 2.105 ;
        RECT 1.305 1.665 1.475 1.910 ;
        RECT 0.940 1.600 1.475 1.665 ;
        RECT 0.905 1.495 1.475 1.600 ;
        RECT 0.905 1.430 1.110 1.495 ;
        RECT 1.645 1.445 2.155 1.690 ;
        RECT 3.655 1.435 4.070 1.745 ;
        RECT 6.150 1.445 6.835 1.735 ;
        RECT 7.010 1.640 7.180 1.935 ;
        RECT 7.815 1.795 7.985 2.635 ;
        RECT 7.010 1.470 7.300 1.640 ;
        RECT 0.905 1.245 1.075 1.430 ;
        RECT 0.540 1.075 1.075 1.245 ;
        RECT 0.905 0.825 1.075 1.075 ;
        RECT 1.245 1.275 1.505 1.325 ;
        RECT 1.245 0.995 1.755 1.275 ;
        RECT 2.685 1.030 3.075 1.360 ;
        RECT 4.720 0.955 5.080 1.275 ;
        RECT 5.250 0.955 5.935 1.125 ;
        RECT 6.105 0.995 6.960 1.275 ;
        RECT 7.130 1.245 7.300 1.470 ;
        RECT 7.130 1.075 7.800 1.245 ;
        RECT 1.925 0.825 2.165 0.935 ;
        RECT 0.905 0.655 2.165 0.825 ;
        RECT 0.180 0.085 0.350 0.565 ;
        RECT 1.020 0.085 1.350 0.465 ;
        RECT 1.535 0.255 2.165 0.655 ;
        RECT 2.415 0.615 3.425 0.785 ;
        RECT 2.415 0.255 2.585 0.615 ;
        RECT 2.755 0.085 3.085 0.445 ;
        RECT 3.255 0.255 3.425 0.615 ;
        RECT 4.195 0.615 5.205 0.785 ;
        RECT 5.420 0.765 5.935 0.955 ;
        RECT 7.130 0.825 7.300 1.075 ;
        RECT 3.695 0.085 4.025 0.490 ;
        RECT 4.195 0.255 4.365 0.615 ;
        RECT 4.535 0.085 4.865 0.445 ;
        RECT 5.035 0.255 5.205 0.615 ;
        RECT 6.380 0.655 7.300 0.825 ;
        RECT 5.540 0.505 5.710 0.595 ;
        RECT 6.380 0.505 6.550 0.655 ;
        RECT 5.540 0.255 6.550 0.505 ;
        RECT 6.780 0.085 7.110 0.445 ;
        RECT 7.895 0.085 8.065 0.565 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 1.985 1.445 2.155 1.615 ;
        RECT 3.845 1.445 4.015 1.615 ;
        RECT 6.605 1.445 6.775 1.615 ;
        RECT 1.525 1.105 1.695 1.275 ;
        RECT 2.905 1.105 3.075 1.275 ;
        RECT 4.765 1.105 4.935 1.275 ;
        RECT 6.145 1.105 6.315 1.275 ;
        RECT 1.985 0.765 2.155 0.935 ;
        RECT 5.685 0.765 5.855 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
      LAYER met1 ;
        RECT 1.925 0.920 2.215 0.965 ;
        RECT 5.625 0.920 5.915 0.965 ;
        RECT 1.925 0.780 5.915 0.920 ;
        RECT 1.925 0.735 2.215 0.780 ;
        RECT 5.625 0.735 5.915 0.780 ;
  END
END sky130_fd_sc_hd__fa_2

#--------EOF---------

MACRO sky130_fd_sc_hd__fa_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fa_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.633000 ;
    PORT
      LAYER met1 ;
        RECT 2.390 1.260 2.680 1.305 ;
        RECT 3.770 1.260 4.060 1.305 ;
        RECT 5.630 1.260 5.920 1.305 ;
        RECT 7.010 1.260 7.300 1.305 ;
        RECT 2.390 1.120 7.300 1.260 ;
        RECT 2.390 1.075 2.680 1.120 ;
        RECT 3.770 1.075 4.060 1.120 ;
        RECT 5.630 1.075 5.920 1.120 ;
        RECT 7.010 1.075 7.300 1.120 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.633000 ;
    PORT
      LAYER met1 ;
        RECT 2.850 1.600 3.140 1.645 ;
        RECT 4.710 1.600 5.000 1.645 ;
        RECT 7.470 1.600 7.760 1.645 ;
        RECT 2.850 1.460 7.760 1.600 ;
        RECT 2.850 1.415 3.140 1.460 ;
        RECT 4.710 1.415 5.000 1.460 ;
        RECT 7.470 1.415 7.760 1.460 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.477000 ;
    PORT
      LAYER li1 ;
        RECT 3.250 1.570 4.340 1.740 ;
        RECT 6.595 1.685 6.845 1.955 ;
        RECT 3.250 1.275 3.420 1.570 ;
        RECT 3.050 1.105 3.420 1.275 ;
        RECT 4.170 1.250 4.340 1.570 ;
        RECT 5.220 1.515 6.845 1.685 ;
        RECT 5.220 1.435 5.580 1.515 ;
        RECT 5.220 1.250 5.390 1.435 ;
        RECT 6.595 1.355 6.845 1.515 ;
        RECT 4.170 0.965 5.390 1.250 ;
    END
  END CIN
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 2.195 1.015 ;
        RECT 7.690 0.785 10.030 1.015 ;
        RECT 0.005 0.105 10.030 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.585 0.845 2.445 ;
        RECT 1.435 1.950 1.645 2.465 ;
        RECT 1.400 1.780 1.645 1.950 ;
        RECT 1.400 1.585 1.570 1.780 ;
        RECT 0.085 1.415 1.570 1.585 ;
        RECT 0.085 0.905 0.435 1.415 ;
        RECT 0.085 0.735 1.525 0.905 ;
        RECT 0.515 0.255 0.845 0.735 ;
        RECT 1.355 0.485 1.525 0.735 ;
        RECT 1.355 0.315 1.685 0.485 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.943000 ;
    PORT
      LAYER li1 ;
        RECT 8.320 1.965 8.490 2.465 ;
        RECT 8.320 1.795 8.570 1.965 ;
        RECT 8.400 1.585 8.570 1.795 ;
        RECT 9.160 1.585 9.490 2.425 ;
        RECT 8.400 1.415 10.035 1.585 ;
        RECT 9.700 0.905 10.035 1.415 ;
        RECT 8.400 0.735 10.035 0.905 ;
        RECT 8.400 0.485 8.650 0.735 ;
        RECT 8.320 0.255 8.650 0.485 ;
        RECT 9.160 0.270 9.490 0.735 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.175 1.795 0.345 2.635 ;
        RECT 1.015 1.795 1.185 2.635 ;
        RECT 1.815 2.275 2.145 2.635 ;
        RECT 2.735 2.080 3.170 2.465 ;
        RECT 2.140 1.910 3.170 2.080 ;
        RECT 3.340 2.105 3.510 2.465 ;
        RECT 3.680 2.275 4.010 2.635 ;
        RECT 4.180 2.105 4.415 2.465 ;
        RECT 3.340 1.935 4.415 2.105 ;
        RECT 4.620 1.915 4.950 2.635 ;
        RECT 5.120 2.105 5.290 2.465 ;
        RECT 5.460 2.275 5.790 2.635 ;
        RECT 5.960 2.105 6.130 2.465 ;
        RECT 6.410 2.125 7.610 2.465 ;
        RECT 7.815 2.275 8.145 2.635 ;
        RECT 5.120 1.935 6.130 2.105 ;
        RECT 7.440 2.105 7.610 2.125 ;
        RECT 7.440 1.935 8.105 2.105 ;
        RECT 2.140 1.665 2.310 1.910 ;
        RECT 1.775 1.600 2.310 1.665 ;
        RECT 1.740 1.495 2.310 1.600 ;
        RECT 1.740 1.430 1.945 1.495 ;
        RECT 2.480 1.445 3.080 1.690 ;
        RECT 4.580 1.435 4.995 1.745 ;
        RECT 7.075 1.445 7.760 1.735 ;
        RECT 7.935 1.640 8.105 1.935 ;
        RECT 8.740 1.795 8.910 2.635 ;
        RECT 9.660 1.795 9.830 2.635 ;
        RECT 7.935 1.470 8.225 1.640 ;
        RECT 1.740 1.245 1.910 1.430 ;
        RECT 0.605 1.075 1.910 1.245 ;
        RECT 1.740 0.825 1.910 1.075 ;
        RECT 2.080 1.275 2.340 1.325 ;
        RECT 2.080 0.995 2.680 1.275 ;
        RECT 3.610 1.030 4.000 1.360 ;
        RECT 5.645 0.955 6.005 1.275 ;
        RECT 6.175 0.955 6.860 1.125 ;
        RECT 7.030 0.995 7.885 1.275 ;
        RECT 8.055 1.245 8.225 1.470 ;
        RECT 8.055 1.075 9.445 1.245 ;
        RECT 2.850 0.825 3.090 0.935 ;
        RECT 1.740 0.655 3.090 0.825 ;
        RECT 0.175 0.085 0.345 0.565 ;
        RECT 1.015 0.085 1.185 0.565 ;
        RECT 1.855 0.085 2.185 0.465 ;
        RECT 2.370 0.255 3.090 0.655 ;
        RECT 3.340 0.615 4.350 0.785 ;
        RECT 3.340 0.255 3.510 0.615 ;
        RECT 3.680 0.085 4.010 0.445 ;
        RECT 4.180 0.255 4.350 0.615 ;
        RECT 5.120 0.615 6.130 0.785 ;
        RECT 6.345 0.765 6.860 0.955 ;
        RECT 8.055 0.825 8.225 1.075 ;
        RECT 4.620 0.085 4.950 0.490 ;
        RECT 5.120 0.255 5.290 0.615 ;
        RECT 5.460 0.085 5.790 0.445 ;
        RECT 5.960 0.255 6.130 0.615 ;
        RECT 7.305 0.655 8.225 0.825 ;
        RECT 6.465 0.505 6.635 0.595 ;
        RECT 7.305 0.505 7.475 0.655 ;
        RECT 6.465 0.255 7.475 0.505 ;
        RECT 7.705 0.085 8.035 0.445 ;
        RECT 8.820 0.085 8.990 0.565 ;
        RECT 9.660 0.085 9.830 0.565 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 2.910 1.445 3.080 1.615 ;
        RECT 4.770 1.445 4.940 1.615 ;
        RECT 7.530 1.445 7.700 1.615 ;
        RECT 2.450 1.105 2.620 1.275 ;
        RECT 3.830 1.105 4.000 1.275 ;
        RECT 5.690 1.105 5.860 1.275 ;
        RECT 7.070 1.105 7.240 1.275 ;
        RECT 2.910 0.765 3.080 0.935 ;
        RECT 6.610 0.765 6.780 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
      LAYER met1 ;
        RECT 2.850 0.920 3.140 0.965 ;
        RECT 6.550 0.920 6.840 0.965 ;
        RECT 2.850 0.780 6.840 0.920 ;
        RECT 2.850 0.735 3.140 0.780 ;
        RECT 6.550 0.735 6.840 0.780 ;
  END
END sky130_fd_sc_hd__fa_4

#--------EOF---------

MACRO sky130_fd_sc_hd__fah_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fah_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.420 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 0.950 1.075 1.440 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.691500 ;
    PORT
      LAYER met1 ;
        RECT 1.930 1.260 2.220 1.305 ;
        RECT 5.620 1.260 5.910 1.305 ;
        RECT 1.930 1.120 5.910 1.260 ;
        RECT 1.930 1.075 2.220 1.120 ;
        RECT 5.620 1.075 5.910 1.120 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 9.475 1.075 9.865 1.325 ;
        RECT 9.690 0.935 9.865 1.075 ;
        RECT 9.690 0.735 10.010 0.935 ;
    END
  END CI
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.420 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.005 3.050 1.015 ;
        RECT 5.095 1.005 12.400 1.015 ;
        RECT 0.005 0.115 12.400 1.005 ;
        RECT 0.005 0.105 5.530 0.115 ;
        RECT 10.960 0.105 12.400 0.115 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.610 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 12.420 2.960 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.435500 ;
    PORT
      LAYER li1 ;
        RECT 10.870 1.495 11.390 2.465 ;
        RECT 10.870 0.825 11.040 1.495 ;
        RECT 10.870 0.270 11.310 0.825 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.506000 ;
    PORT
      LAYER li1 ;
        RECT 11.985 1.785 12.335 2.465 ;
        RECT 12.110 0.825 12.335 1.785 ;
        RECT 11.980 0.255 12.335 0.825 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 12.420 2.805 ;
        RECT 0.085 2.065 0.395 2.465 ;
        RECT 0.565 2.260 0.930 2.635 ;
        RECT 2.065 2.235 2.395 2.635 ;
        RECT 2.635 2.295 4.950 2.465 ;
        RECT 5.125 2.295 7.560 2.465 ;
        RECT 2.635 2.065 2.805 2.295 ;
        RECT 0.085 1.895 2.805 2.065 ;
        RECT 3.030 1.955 4.320 2.125 ;
        RECT 0.085 1.500 0.445 1.895 ;
        RECT 0.985 1.615 1.315 1.715 ;
        RECT 0.085 0.805 0.255 1.500 ;
        RECT 0.615 1.455 1.315 1.615 ;
        RECT 0.610 1.445 1.315 1.455 ;
        RECT 1.490 1.500 1.840 1.725 ;
        RECT 1.490 1.445 1.820 1.500 ;
        RECT 0.610 1.380 0.815 1.445 ;
        RECT 0.610 1.325 0.780 1.380 ;
        RECT 0.425 0.995 0.780 1.325 ;
        RECT 0.595 0.905 0.780 0.995 ;
        RECT 1.615 0.905 1.820 1.445 ;
        RECT 2.015 1.410 2.190 1.725 ;
        RECT 2.360 1.445 2.860 1.715 ;
        RECT 1.990 1.275 2.190 1.410 ;
        RECT 1.990 1.075 2.495 1.275 ;
        RECT 0.085 0.255 0.425 0.805 ;
        RECT 0.595 0.735 1.320 0.905 ;
        RECT 0.595 0.085 0.765 0.545 ;
        RECT 0.990 0.255 1.320 0.735 ;
        RECT 1.500 0.885 1.820 0.905 ;
        RECT 1.500 0.715 2.520 0.885 ;
        RECT 1.500 0.255 1.840 0.715 ;
        RECT 2.010 0.085 2.180 0.545 ;
        RECT 2.350 0.425 2.520 0.715 ;
        RECT 2.690 0.595 2.860 1.445 ;
        RECT 3.030 0.465 3.200 1.955 ;
        RECT 3.985 1.785 4.320 1.955 ;
        RECT 3.370 1.455 3.815 1.785 ;
        RECT 3.370 0.805 3.540 1.455 ;
        RECT 4.070 1.160 4.535 1.615 ;
        RECT 4.070 1.075 4.400 1.160 ;
        RECT 4.705 0.925 4.875 2.295 ;
        RECT 5.125 1.320 5.295 2.295 ;
        RECT 5.475 1.700 5.875 2.030 ;
        RECT 6.290 1.955 7.220 2.125 ;
        RECT 6.290 1.615 6.460 1.955 ;
        RECT 6.105 1.445 6.460 1.615 ;
        RECT 5.125 1.150 5.505 1.320 ;
        RECT 5.320 0.925 5.505 1.150 ;
        RECT 5.675 0.995 5.925 1.325 ;
        RECT 6.710 1.275 6.880 1.785 ;
        RECT 4.480 0.905 5.145 0.925 ;
        RECT 4.070 0.805 5.145 0.905 ;
        RECT 5.320 0.865 5.520 0.925 ;
        RECT 5.335 0.840 5.520 0.865 ;
        RECT 3.370 0.635 3.900 0.805 ;
        RECT 4.070 0.780 5.155 0.805 ;
        RECT 4.070 0.755 5.170 0.780 ;
        RECT 4.070 0.735 4.560 0.755 ;
        RECT 4.925 0.740 5.170 0.755 ;
        RECT 4.925 0.735 5.180 0.740 ;
        RECT 4.070 0.645 4.400 0.735 ;
        RECT 4.950 0.715 5.180 0.735 ;
        RECT 4.980 0.690 5.180 0.715 ;
        RECT 5.000 0.655 5.180 0.690 ;
        RECT 4.650 0.465 4.840 0.585 ;
        RECT 3.030 0.425 4.840 0.465 ;
        RECT 2.350 0.255 4.840 0.425 ;
        RECT 5.010 0.425 5.180 0.655 ;
        RECT 5.350 0.595 5.520 0.840 ;
        RECT 6.105 0.740 6.435 1.275 ;
        RECT 6.610 0.925 6.880 1.275 ;
        RECT 7.050 1.175 7.220 1.955 ;
        RECT 7.390 1.425 7.560 2.295 ;
        RECT 7.730 2.295 9.655 2.465 ;
        RECT 7.730 1.510 7.960 2.295 ;
        RECT 8.145 1.955 9.250 2.125 ;
        RECT 7.390 1.400 7.575 1.425 ;
        RECT 7.390 1.375 7.595 1.400 ;
        RECT 7.390 1.275 7.620 1.375 ;
        RECT 7.050 1.130 7.245 1.175 ;
        RECT 7.050 1.060 7.280 1.130 ;
        RECT 7.065 1.045 7.280 1.060 ;
        RECT 7.090 1.010 7.280 1.045 ;
        RECT 6.610 0.755 6.940 0.925 ;
        RECT 6.770 0.595 6.940 0.755 ;
        RECT 7.110 0.765 7.280 1.010 ;
        RECT 7.450 0.995 7.620 1.275 ;
        RECT 7.790 0.825 7.960 1.510 ;
        RECT 8.225 1.445 8.910 1.785 ;
        RECT 8.225 0.925 8.405 1.445 ;
        RECT 9.080 1.275 9.250 1.955 ;
        RECT 9.420 1.705 9.655 2.295 ;
        RECT 9.840 2.275 10.175 2.635 ;
        RECT 10.345 1.875 10.690 2.465 ;
        RECT 9.420 1.495 10.350 1.705 ;
        RECT 7.110 0.595 7.445 0.765 ;
        RECT 5.750 0.425 6.100 0.565 ;
        RECT 5.010 0.255 6.100 0.425 ;
        RECT 6.270 0.425 6.600 0.570 ;
        RECT 7.705 0.425 7.960 0.825 ;
        RECT 8.155 0.595 8.405 0.925 ;
        RECT 8.575 1.105 9.250 1.275 ;
        RECT 8.575 0.595 8.745 1.105 ;
        RECT 10.180 0.995 10.350 1.495 ;
        RECT 8.920 0.685 9.300 0.935 ;
        RECT 10.520 0.825 10.690 1.875 ;
        RECT 11.560 1.785 11.815 2.635 ;
        RECT 11.210 0.995 11.460 1.325 ;
        RECT 11.630 0.995 11.940 1.615 ;
        RECT 9.400 0.425 9.735 0.515 ;
        RECT 6.270 0.255 9.735 0.425 ;
        RECT 9.905 0.085 10.075 0.565 ;
        RECT 10.245 0.285 10.690 0.825 ;
        RECT 11.480 0.085 11.810 0.825 ;
        RECT 0.000 -0.085 12.420 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 2.450 1.445 2.620 1.615 ;
        RECT 1.990 1.105 2.160 1.275 ;
        RECT 4.365 1.445 4.535 1.615 ;
        RECT 3.370 0.765 3.540 0.935 ;
        RECT 5.570 1.785 5.740 1.955 ;
        RECT 6.150 1.445 6.320 1.615 ;
        RECT 5.680 1.105 5.850 1.275 ;
        RECT 6.150 0.765 6.320 0.935 ;
        RECT 6.610 1.105 6.780 1.275 ;
        RECT 9.080 1.785 9.250 1.955 ;
        RECT 8.460 1.445 8.630 1.615 ;
        RECT 10.520 1.785 10.690 1.955 ;
        RECT 8.920 0.765 9.090 0.935 ;
        RECT 11.680 1.445 11.850 1.615 ;
        RECT 11.220 1.105 11.390 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
      LAYER met1 ;
        RECT 3.925 1.940 4.215 1.985 ;
        RECT 5.510 1.940 5.800 1.985 ;
        RECT 3.925 1.800 5.800 1.940 ;
        RECT 3.925 1.755 4.215 1.800 ;
        RECT 5.510 1.755 5.800 1.800 ;
        RECT 9.020 1.940 9.310 1.985 ;
        RECT 10.460 1.940 10.750 1.985 ;
        RECT 9.020 1.800 10.750 1.940 ;
        RECT 9.020 1.755 9.310 1.800 ;
        RECT 10.460 1.755 10.750 1.800 ;
        RECT 2.390 1.600 2.680 1.645 ;
        RECT 4.305 1.600 4.595 1.645 ;
        RECT 6.090 1.600 6.380 1.645 ;
        RECT 2.390 1.460 6.380 1.600 ;
        RECT 2.390 1.415 2.680 1.460 ;
        RECT 4.305 1.415 4.595 1.460 ;
        RECT 6.090 1.415 6.380 1.460 ;
        RECT 8.400 1.600 8.690 1.645 ;
        RECT 11.620 1.600 11.910 1.645 ;
        RECT 8.400 1.460 11.910 1.600 ;
        RECT 8.400 1.415 8.690 1.460 ;
        RECT 11.620 1.415 11.910 1.460 ;
        RECT 6.550 1.260 6.840 1.305 ;
        RECT 11.160 1.260 11.450 1.305 ;
        RECT 6.550 1.120 11.450 1.260 ;
        RECT 6.550 1.075 6.840 1.120 ;
        RECT 11.160 1.075 11.450 1.120 ;
        RECT 3.310 0.920 3.600 0.965 ;
        RECT 6.090 0.920 6.380 0.965 ;
        RECT 8.860 0.920 9.150 0.965 ;
        RECT 3.310 0.780 9.150 0.920 ;
        RECT 3.310 0.735 3.600 0.780 ;
        RECT 6.090 0.735 6.380 0.780 ;
        RECT 8.860 0.735 9.150 0.780 ;
  END
END sky130_fd_sc_hd__fah_1

#--------EOF---------

MACRO sky130_fd_sc_hd__fahcin_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fahcin_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.420 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.950 1.075 1.340 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.691500 ;
    PORT
      LAYER met1 ;
        RECT 1.465 0.920 1.755 0.965 ;
        RECT 4.225 0.920 4.515 0.965 ;
        RECT 1.465 0.780 4.515 0.920 ;
        RECT 1.465 0.735 1.755 0.780 ;
        RECT 4.225 0.735 4.515 0.780 ;
    END
  END B
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.493500 ;
    PORT
      LAYER li1 ;
        RECT 10.520 1.075 10.965 1.275 ;
    END
  END CIN
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.420 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.495 1.005 12.415 1.015 ;
        RECT 0.005 0.115 12.415 1.005 ;
        RECT 0.005 0.105 1.720 0.115 ;
        RECT 3.050 0.105 5.580 0.115 ;
        RECT 10.055 0.105 12.415 0.115 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.610 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 12.420 2.960 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.402800 ;
    PORT
      LAYER li1 ;
        RECT 6.700 1.675 6.870 1.785 ;
        RECT 6.600 0.925 6.870 1.675 ;
        RECT 6.600 0.755 6.925 0.925 ;
        RECT 6.755 0.595 6.925 0.755 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.470250 ;
    PORT
      LAYER li1 ;
        RECT 12.000 1.785 12.335 2.465 ;
        RECT 12.125 0.825 12.335 1.785 ;
        RECT 11.995 0.255 12.335 0.825 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 12.420 2.805 ;
        RECT 0.085 2.010 0.430 2.465 ;
        RECT 0.600 2.180 0.770 2.635 ;
        RECT 1.715 2.385 3.515 2.465 ;
        RECT 0.940 2.295 3.515 2.385 ;
        RECT 0.940 2.215 1.970 2.295 ;
        RECT 0.940 2.010 1.110 2.215 ;
        RECT 3.245 2.110 3.460 2.295 ;
        RECT 0.085 1.840 1.110 2.010 ;
        RECT 1.280 1.955 1.450 2.045 ;
        RECT 0.085 1.500 0.440 1.840 ;
        RECT 1.280 1.785 2.050 1.955 ;
        RECT 2.565 1.785 2.895 2.045 ;
        RECT 1.280 1.670 1.450 1.785 ;
        RECT 0.610 1.500 1.450 1.670 ;
        RECT 0.085 0.805 0.255 1.500 ;
        RECT 0.610 1.325 0.780 1.500 ;
        RECT 2.220 1.350 2.390 1.785 ;
        RECT 0.425 0.995 0.780 1.325 ;
        RECT 0.610 0.905 0.780 0.995 ;
        RECT 0.085 0.735 0.430 0.805 ;
        RECT 0.610 0.735 1.325 0.905 ;
        RECT 0.100 0.255 0.430 0.735 ;
        RECT 0.630 0.085 0.800 0.545 ;
        RECT 0.995 0.465 1.325 0.735 ;
        RECT 1.510 0.665 1.740 1.325 ;
        RECT 1.985 0.675 2.390 1.350 ;
        RECT 2.950 1.265 3.120 1.615 ;
        RECT 2.800 1.245 3.120 1.265 ;
        RECT 2.640 1.095 3.120 1.245 ;
        RECT 2.640 1.075 2.970 1.095 ;
        RECT 3.290 0.925 3.460 2.110 ;
        RECT 3.710 2.290 5.065 2.460 ;
        RECT 3.710 1.320 3.880 2.290 ;
        RECT 4.080 1.695 4.445 2.120 ;
        RECT 4.815 2.065 5.065 2.290 ;
        RECT 5.260 2.235 5.590 2.635 ;
        RECT 5.825 2.295 7.950 2.465 ;
        RECT 5.825 2.065 5.995 2.295 ;
        RECT 4.815 1.895 5.995 2.065 ;
        RECT 6.200 1.955 7.210 2.125 ;
        RECT 6.200 1.895 6.530 1.955 ;
        RECT 6.200 1.725 6.370 1.895 ;
        RECT 4.690 1.385 5.170 1.725 ;
        RECT 5.635 1.555 6.370 1.725 ;
        RECT 4.830 1.325 5.170 1.385 ;
        RECT 3.710 1.150 4.070 1.320 ;
        RECT 3.055 0.905 3.730 0.925 ;
        RECT 2.220 0.595 2.390 0.675 ;
        RECT 2.620 0.755 3.730 0.905 ;
        RECT 2.620 0.735 3.135 0.755 ;
        RECT 2.620 0.655 3.025 0.735 ;
        RECT 3.215 0.465 3.390 0.585 ;
        RECT 0.995 0.425 2.100 0.465 ;
        RECT 2.515 0.425 3.390 0.465 ;
        RECT 0.995 0.255 3.390 0.425 ;
        RECT 3.560 0.425 3.730 0.755 ;
        RECT 3.900 0.595 4.070 1.150 ;
        RECT 4.240 0.645 4.490 1.325 ;
        RECT 4.830 0.995 5.630 1.325 ;
        RECT 4.830 0.510 5.000 0.995 ;
        RECT 5.800 0.815 5.970 1.555 ;
        RECT 4.240 0.425 4.570 0.475 ;
        RECT 3.560 0.255 4.570 0.425 ;
        RECT 5.180 0.085 5.510 0.805 ;
        RECT 5.680 0.380 5.970 0.815 ;
        RECT 6.140 0.740 6.425 1.325 ;
        RECT 7.040 1.230 7.210 1.955 ;
        RECT 7.380 1.530 7.550 2.125 ;
        RECT 7.780 1.720 7.950 2.295 ;
        RECT 8.220 2.295 9.410 2.465 ;
        RECT 8.220 1.955 8.390 2.295 ;
        RECT 8.560 1.785 8.890 2.125 ;
        RECT 7.780 1.550 8.035 1.720 ;
        RECT 7.380 1.360 7.610 1.530 ;
        RECT 7.440 1.290 7.610 1.360 ;
        RECT 7.040 1.060 7.270 1.230 ;
        RECT 7.440 1.105 7.695 1.290 ;
        RECT 7.100 0.925 7.270 1.060 ;
        RECT 7.100 0.595 7.350 0.925 ;
        RECT 6.255 0.425 6.585 0.570 ;
        RECT 7.520 0.425 7.695 1.105 ;
        RECT 7.865 0.995 8.035 1.550 ;
        RECT 8.375 1.530 8.890 1.785 ;
        RECT 9.240 2.045 9.410 2.295 ;
        RECT 10.190 2.195 10.360 2.635 ;
        RECT 9.240 2.040 10.105 2.045 ;
        RECT 9.240 2.035 10.120 2.040 ;
        RECT 9.240 2.030 10.130 2.035 ;
        RECT 9.240 2.025 10.145 2.030 ;
        RECT 10.535 2.025 10.885 2.465 ;
        RECT 9.240 1.875 10.885 2.025 ;
        RECT 8.375 1.445 8.670 1.530 ;
        RECT 8.375 0.925 8.555 1.445 ;
        RECT 8.835 0.995 9.070 1.325 ;
        RECT 6.255 0.255 7.695 0.425 ;
        RECT 7.865 0.425 8.035 0.740 ;
        RECT 8.305 0.595 8.555 0.925 ;
        RECT 9.240 0.765 9.410 1.875 ;
        RECT 10.055 1.870 10.885 1.875 ;
        RECT 10.070 1.865 10.885 1.870 ;
        RECT 10.085 1.860 10.885 1.865 ;
        RECT 10.100 1.855 10.885 1.860 ;
        RECT 8.725 0.595 9.410 0.765 ;
        RECT 9.640 1.535 10.010 1.705 ;
        RECT 9.640 0.825 9.810 1.535 ;
        RECT 10.180 1.445 10.885 1.855 ;
        RECT 11.075 1.455 11.405 2.465 ;
        RECT 11.575 1.785 11.830 2.635 ;
        RECT 10.180 1.325 10.350 1.445 ;
        RECT 9.980 0.995 10.350 1.325 ;
        RECT 10.180 0.905 10.350 0.995 ;
        RECT 9.640 0.425 9.980 0.825 ;
        RECT 10.180 0.735 10.910 0.905 ;
        RECT 7.865 0.255 9.980 0.425 ;
        RECT 10.180 0.085 10.350 0.565 ;
        RECT 10.530 0.285 10.910 0.735 ;
        RECT 11.155 0.680 11.405 1.455 ;
        RECT 11.645 0.995 11.955 1.615 ;
        RECT 11.155 0.270 11.325 0.680 ;
        RECT 11.495 0.085 11.825 0.510 ;
        RECT 0.000 -0.085 12.420 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 1.880 1.785 2.050 1.955 ;
        RECT 2.570 1.785 2.740 1.955 ;
        RECT 1.525 0.765 1.695 0.935 ;
        RECT 1.985 1.105 2.155 1.275 ;
        RECT 2.950 1.445 3.120 1.615 ;
        RECT 4.140 1.785 4.310 1.955 ;
        RECT 4.760 1.445 4.930 1.615 ;
        RECT 4.285 0.765 4.455 0.935 ;
        RECT 6.140 1.105 6.310 1.275 ;
        RECT 8.440 1.445 8.610 1.615 ;
        RECT 7.520 0.765 7.690 0.935 ;
        RECT 8.900 1.105 9.070 1.275 ;
        RECT 11.680 1.445 11.850 1.615 ;
        RECT 11.220 0.765 11.390 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
      LAYER met1 ;
        RECT 1.820 1.940 2.110 1.985 ;
        RECT 2.510 1.940 2.800 1.985 ;
        RECT 4.080 1.940 4.370 1.985 ;
        RECT 1.820 1.800 4.370 1.940 ;
        RECT 1.820 1.755 2.110 1.800 ;
        RECT 2.510 1.755 2.800 1.800 ;
        RECT 4.080 1.755 4.370 1.800 ;
        RECT 2.890 1.600 3.180 1.645 ;
        RECT 4.700 1.600 4.990 1.645 ;
        RECT 2.890 1.460 4.990 1.600 ;
        RECT 2.890 1.415 3.180 1.460 ;
        RECT 4.700 1.415 4.990 1.460 ;
        RECT 8.380 1.600 8.670 1.645 ;
        RECT 11.620 1.600 11.910 1.645 ;
        RECT 8.380 1.460 11.910 1.600 ;
        RECT 8.380 1.415 8.670 1.460 ;
        RECT 11.620 1.415 11.910 1.460 ;
        RECT 1.925 1.260 2.215 1.305 ;
        RECT 6.080 1.260 6.370 1.305 ;
        RECT 8.840 1.260 9.130 1.305 ;
        RECT 1.925 1.120 9.130 1.260 ;
        RECT 1.925 1.075 2.215 1.120 ;
        RECT 6.080 1.075 6.370 1.120 ;
        RECT 8.840 1.075 9.130 1.120 ;
        RECT 7.460 0.920 7.750 0.965 ;
        RECT 11.160 0.920 11.450 0.965 ;
        RECT 7.460 0.780 11.450 0.920 ;
        RECT 7.460 0.735 7.750 0.780 ;
        RECT 11.160 0.735 11.450 0.780 ;
  END
END sky130_fd_sc_hd__fahcin_1

#--------EOF---------

MACRO sky130_fd_sc_hd__fahcon_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__fahcon_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.420 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.950 1.075 1.340 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.937500 ;
    PORT
      LAYER met1 ;
        RECT 1.465 0.920 1.755 0.965 ;
        RECT 4.250 0.920 4.540 0.965 ;
        RECT 1.465 0.780 4.540 0.920 ;
        RECT 1.465 0.735 1.755 0.780 ;
        RECT 4.250 0.735 4.540 0.780 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.493500 ;
    PORT
      LAYER li1 ;
        RECT 10.530 1.075 10.975 1.275 ;
    END
  END CI
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.420 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.495 1.005 12.415 1.015 ;
        RECT 0.010 0.115 12.415 1.005 ;
        RECT 0.010 0.105 1.720 0.115 ;
        RECT 3.070 0.105 5.610 0.115 ;
        RECT 10.065 0.105 12.415 0.115 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.610 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 12.420 2.960 ;
    END
  END VPWR
  PIN COUT_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.402800 ;
    PORT
      LAYER li1 ;
        RECT 6.710 1.675 6.880 1.785 ;
        RECT 6.610 0.925 6.880 1.675 ;
        RECT 6.610 0.755 6.935 0.925 ;
        RECT 6.765 0.595 6.935 0.755 ;
    END
  END COUT_N
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.463750 ;
    PORT
      LAYER li1 ;
        RECT 12.010 1.785 12.335 2.465 ;
        RECT 12.135 0.825 12.335 1.785 ;
        RECT 11.995 0.255 12.335 0.825 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 12.420 2.805 ;
        RECT 0.085 2.010 0.430 2.465 ;
        RECT 0.600 2.180 0.770 2.635 ;
        RECT 2.375 2.385 3.540 2.465 ;
        RECT 0.940 2.295 3.540 2.385 ;
        RECT 3.725 2.295 5.100 2.465 ;
        RECT 0.940 2.215 2.545 2.295 ;
        RECT 0.940 2.010 1.110 2.215 ;
        RECT 0.085 1.840 1.110 2.010 ;
        RECT 1.280 1.875 2.920 2.045 ;
        RECT 0.085 1.500 0.440 1.840 ;
        RECT 1.280 1.670 1.450 1.875 ;
        RECT 0.610 1.500 1.450 1.670 ;
        RECT 0.085 0.805 0.255 1.500 ;
        RECT 0.610 1.325 0.780 1.500 ;
        RECT 0.425 0.995 0.780 1.325 ;
        RECT 0.610 0.905 0.780 0.995 ;
        RECT 0.085 0.735 0.430 0.805 ;
        RECT 0.610 0.735 1.325 0.905 ;
        RECT 0.100 0.255 0.430 0.735 ;
        RECT 0.630 0.085 0.800 0.545 ;
        RECT 0.995 0.465 1.325 0.735 ;
        RECT 1.510 0.710 1.780 1.325 ;
        RECT 1.965 0.635 2.470 1.705 ;
        RECT 2.640 1.160 3.100 1.615 ;
        RECT 2.640 1.075 2.975 1.160 ;
        RECT 3.270 0.925 3.440 2.295 ;
        RECT 3.725 1.320 3.895 2.295 ;
        RECT 4.210 1.755 4.380 2.095 ;
        RECT 4.875 2.065 5.100 2.295 ;
        RECT 5.270 2.235 5.600 2.635 ;
        RECT 5.835 2.295 7.960 2.465 ;
        RECT 5.835 2.065 6.005 2.295 ;
        RECT 4.875 1.895 6.005 2.065 ;
        RECT 6.210 1.955 7.220 2.125 ;
        RECT 6.210 1.895 6.540 1.955 ;
        RECT 6.210 1.725 6.380 1.895 ;
        RECT 4.700 1.385 5.180 1.725 ;
        RECT 5.645 1.555 6.380 1.725 ;
        RECT 3.725 1.150 4.095 1.320 ;
        RECT 3.055 0.905 3.750 0.925 ;
        RECT 2.640 0.755 3.750 0.905 ;
        RECT 2.640 0.735 3.160 0.755 ;
        RECT 2.640 0.655 3.025 0.735 ;
        RECT 3.240 0.465 3.410 0.585 ;
        RECT 0.995 0.255 3.410 0.465 ;
        RECT 3.580 0.425 3.750 0.755 ;
        RECT 3.925 0.595 4.095 1.150 ;
        RECT 4.265 0.645 4.515 1.325 ;
        RECT 4.840 0.995 5.180 1.385 ;
        RECT 4.840 0.510 5.030 0.995 ;
        RECT 5.810 0.815 5.980 1.555 ;
        RECT 4.265 0.425 4.595 0.475 ;
        RECT 3.580 0.255 4.595 0.425 ;
        RECT 5.200 0.085 5.530 0.805 ;
        RECT 5.700 0.380 5.980 0.815 ;
        RECT 6.150 0.740 6.435 1.325 ;
        RECT 7.050 1.230 7.220 1.955 ;
        RECT 7.390 1.530 7.560 2.125 ;
        RECT 7.790 1.720 7.960 2.295 ;
        RECT 8.230 2.295 9.950 2.465 ;
        RECT 8.230 1.785 8.400 2.295 ;
        RECT 9.620 2.215 9.950 2.295 ;
        RECT 10.120 2.275 10.455 2.635 ;
        RECT 7.790 1.550 8.045 1.720 ;
        RECT 8.570 1.615 8.900 2.125 ;
        RECT 7.390 1.360 7.620 1.530 ;
        RECT 7.450 1.290 7.620 1.360 ;
        RECT 7.050 1.060 7.280 1.230 ;
        RECT 7.450 1.105 7.700 1.290 ;
        RECT 7.110 0.925 7.280 1.060 ;
        RECT 7.110 0.595 7.360 0.925 ;
        RECT 6.265 0.425 6.595 0.570 ;
        RECT 7.530 0.425 7.700 1.105 ;
        RECT 7.875 0.995 8.045 1.550 ;
        RECT 8.440 1.530 8.900 1.615 ;
        RECT 9.070 2.045 9.420 2.125 ;
        RECT 9.070 1.530 9.450 2.045 ;
        RECT 8.440 1.445 8.740 1.530 ;
        RECT 6.265 0.255 7.700 0.425 ;
        RECT 7.935 0.425 8.270 0.825 ;
        RECT 8.440 0.765 8.610 1.445 ;
        RECT 8.780 0.995 9.110 1.275 ;
        RECT 8.440 0.595 8.900 0.765 ;
        RECT 9.280 0.425 9.450 1.530 ;
        RECT 7.935 0.255 9.450 0.425 ;
        RECT 9.650 1.535 9.950 2.215 ;
        RECT 10.625 2.045 10.835 2.465 ;
        RECT 9.650 0.825 9.820 1.535 ;
        RECT 10.190 1.455 10.835 2.045 ;
        RECT 11.085 1.455 11.415 2.465 ;
        RECT 11.585 1.785 11.840 2.635 ;
        RECT 10.190 1.325 10.360 1.455 ;
        RECT 9.990 0.995 10.360 1.325 ;
        RECT 10.190 0.905 10.360 0.995 ;
        RECT 9.650 0.255 10.020 0.825 ;
        RECT 10.190 0.735 10.920 0.905 ;
        RECT 10.200 0.085 10.370 0.565 ;
        RECT 10.540 0.285 10.920 0.735 ;
        RECT 11.165 0.680 11.415 1.455 ;
        RECT 11.655 0.995 11.965 1.615 ;
        RECT 11.165 0.270 11.335 0.680 ;
        RECT 11.535 0.085 11.825 0.555 ;
        RECT 0.000 -0.085 12.420 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 1.280 1.785 1.450 1.955 ;
        RECT 1.525 0.765 1.695 0.935 ;
        RECT 1.985 1.105 2.155 1.275 ;
        RECT 2.930 1.445 3.100 1.615 ;
        RECT 4.210 1.785 4.380 1.955 ;
        RECT 4.770 1.445 4.940 1.615 ;
        RECT 4.310 0.765 4.480 0.935 ;
        RECT 6.150 1.105 6.320 1.275 ;
        RECT 8.450 1.445 8.620 1.615 ;
        RECT 9.280 1.785 9.450 1.955 ;
        RECT 7.530 0.765 7.700 0.935 ;
        RECT 8.910 1.105 9.080 1.275 ;
        RECT 10.190 1.785 10.360 1.955 ;
        RECT 11.690 1.445 11.860 1.615 ;
        RECT 11.230 0.765 11.400 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
      LAYER met1 ;
        RECT 1.195 1.940 1.510 1.985 ;
        RECT 4.150 1.940 4.440 1.985 ;
        RECT 1.195 1.800 4.440 1.940 ;
        RECT 1.195 1.755 1.510 1.800 ;
        RECT 4.150 1.755 4.440 1.800 ;
        RECT 9.195 1.940 9.510 1.985 ;
        RECT 10.130 1.940 10.420 1.985 ;
        RECT 9.195 1.800 10.420 1.940 ;
        RECT 9.195 1.755 9.510 1.800 ;
        RECT 10.130 1.755 10.420 1.800 ;
        RECT 2.845 1.600 3.160 1.645 ;
        RECT 4.710 1.600 5.000 1.645 ;
        RECT 2.845 1.460 5.000 1.600 ;
        RECT 2.845 1.415 3.160 1.460 ;
        RECT 4.710 1.415 5.000 1.460 ;
        RECT 8.390 1.600 8.680 1.645 ;
        RECT 11.630 1.600 11.920 1.645 ;
        RECT 8.390 1.460 11.920 1.600 ;
        RECT 8.390 1.415 8.680 1.460 ;
        RECT 11.630 1.415 11.920 1.460 ;
        RECT 1.925 1.260 2.215 1.305 ;
        RECT 6.090 1.260 6.380 1.305 ;
        RECT 8.850 1.260 9.140 1.305 ;
        RECT 1.925 1.120 9.140 1.260 ;
        RECT 1.925 1.075 2.215 1.120 ;
        RECT 6.090 1.075 6.380 1.120 ;
        RECT 8.850 1.075 9.140 1.120 ;
        RECT 7.470 0.920 7.760 0.965 ;
        RECT 11.170 0.920 11.460 0.965 ;
        RECT 7.470 0.780 11.460 0.920 ;
        RECT 7.470 0.735 7.760 0.780 ;
        RECT 11.170 0.735 11.460 0.780 ;
  END
END sky130_fd_sc_hd__fahcon_1

#--------EOF---------

MACRO sky130_fd_sc_hd__fill_1
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.140 -0.055 0.260 0.055 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.460 2.805 ;
        RECT 0.000 -0.085 0.460 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
  END
END sky130_fd_sc_hd__fill_1

#--------EOF---------

MACRO sky130_fd_sc_hd__fill_2
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.920 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 0.920 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155 -0.050 0.315 0.060 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.110 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.920 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.920 2.805 ;
        RECT 0.000 -0.085 0.920 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
  END
END sky130_fd_sc_hd__fill_2

#--------EOF---------

MACRO sky130_fd_sc_hd__fill_4
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.175 -0.060 0.285 0.060 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__fill_4

#--------EOF---------

MACRO sky130_fd_sc_hd__fill_8
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.130 -0.120 0.350 0.050 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__fill_8

#--------EOF---------

MACRO sky130_fd_sc_hd__ha_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ha_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT 3.360 1.485 3.585 1.615 ;
        RECT 2.335 1.315 3.585 1.485 ;
        RECT 3.360 1.055 3.585 1.315 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT 1.850 1.825 2.155 2.375 ;
        RECT 1.850 1.655 3.165 1.825 ;
        RECT 1.850 1.345 2.155 1.655 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 0.935 1.015 ;
        RECT 3.675 0.785 4.595 1.015 ;
        RECT 0.005 0.105 4.595 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 4.175 1.565 4.515 2.415 ;
        RECT 4.330 0.825 4.515 1.565 ;
        RECT 4.175 0.315 4.515 0.825 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.565 0.425 2.415 ;
        RECT 0.090 0.825 0.320 1.565 ;
        RECT 0.090 0.315 0.425 0.825 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.595 2.275 1.260 2.635 ;
        RECT 0.595 1.515 0.790 2.275 ;
        RECT 1.510 2.105 1.680 2.355 ;
        RECT 2.450 2.275 3.120 2.635 ;
        RECT 0.960 1.935 1.680 2.105 ;
        RECT 3.350 1.955 3.520 2.355 ;
        RECT 3.755 2.125 4.005 2.635 ;
        RECT 0.960 1.245 1.130 1.935 ;
        RECT 3.350 1.785 4.005 1.955 ;
        RECT 3.835 1.325 4.005 1.785 ;
        RECT 0.490 1.075 1.130 1.245 ;
        RECT 0.595 0.085 0.790 0.885 ;
        RECT 0.960 0.675 1.130 1.075 ;
        RECT 1.300 1.145 1.470 1.325 ;
        RECT 1.300 0.975 3.170 1.145 ;
        RECT 3.000 0.885 3.170 0.975 ;
        RECT 3.835 0.995 4.160 1.325 ;
        RECT 3.835 0.885 4.005 0.995 ;
        RECT 0.960 0.345 1.285 0.675 ;
        RECT 1.535 0.635 2.545 0.805 ;
        RECT 1.535 0.345 1.705 0.635 ;
        RECT 1.875 0.085 2.205 0.465 ;
        RECT 2.375 0.345 2.545 0.635 ;
        RECT 3.000 0.715 4.005 0.885 ;
        RECT 3.000 0.345 3.170 0.715 ;
        RECT 3.755 0.085 4.005 0.545 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__ha_1

#--------EOF---------

MACRO sky130_fd_sc_hd__ha_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ha_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 3.820 1.225 4.045 1.675 ;
        RECT 2.790 1.055 4.045 1.225 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 2.310 1.395 3.595 1.675 ;
        RECT 2.310 1.005 2.615 1.395 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 1.395 1.015 ;
        RECT 4.135 0.785 5.515 1.015 ;
        RECT 0.005 0.105 5.515 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.511500 ;
    PORT
      LAYER li1 ;
        RECT 4.715 1.545 4.965 2.415 ;
        RECT 4.790 0.825 4.965 1.545 ;
        RECT 4.635 0.315 4.965 0.825 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.511500 ;
    PORT
      LAYER li1 ;
        RECT 0.555 1.565 0.885 2.415 ;
        RECT 0.555 0.825 0.780 1.565 ;
        RECT 0.555 0.315 0.885 0.825 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.135 1.495 0.375 2.635 ;
        RECT 1.055 1.515 1.250 2.635 ;
        RECT 1.420 2.205 2.220 2.375 ;
        RECT 2.850 2.205 3.640 2.635 ;
        RECT 1.420 1.245 1.590 2.205 ;
        RECT 3.810 2.025 3.980 2.355 ;
        RECT 4.215 2.205 4.545 2.635 ;
        RECT 0.950 1.075 1.590 1.245 ;
        RECT 0.135 0.085 0.375 0.885 ;
        RECT 1.055 0.085 1.250 0.885 ;
        RECT 1.420 0.675 1.590 1.075 ;
        RECT 1.760 1.855 4.465 2.025 ;
        RECT 1.760 0.995 1.930 1.855 ;
        RECT 4.295 1.325 4.465 1.855 ;
        RECT 5.145 1.495 5.385 2.635 ;
        RECT 4.295 0.995 4.620 1.325 ;
        RECT 4.295 0.885 4.465 0.995 ;
        RECT 1.420 0.345 1.745 0.675 ;
        RECT 1.995 0.635 3.005 0.805 ;
        RECT 1.995 0.345 2.165 0.635 ;
        RECT 2.335 0.085 2.665 0.465 ;
        RECT 2.835 0.345 3.005 0.635 ;
        RECT 3.460 0.715 4.465 0.885 ;
        RECT 3.460 0.345 3.630 0.715 ;
        RECT 4.215 0.085 4.465 0.545 ;
        RECT 5.145 0.085 5.385 0.885 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__ha_2

#--------EOF---------

MACRO sky130_fd_sc_hd__ha_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__ha_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 4.210 1.505 6.810 1.675 ;
        RECT 4.210 1.245 4.380 1.505 ;
        RECT 3.320 1.075 4.380 1.245 ;
        RECT 5.625 0.995 5.795 1.505 ;
        RECT 6.580 1.325 6.810 1.505 ;
        RECT 6.580 0.995 7.055 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 4.550 1.165 4.720 1.325 ;
        RECT 4.550 0.995 5.455 1.165 ;
        RECT 5.285 0.875 5.455 0.995 ;
        RECT 5.285 0.845 5.495 0.875 ;
        RECT 5.285 0.825 5.535 0.845 ;
        RECT 6.085 0.825 6.315 1.325 ;
        RECT 5.285 0.730 6.315 0.825 ;
        RECT 5.295 0.720 6.315 0.730 ;
        RECT 5.310 0.710 6.315 0.720 ;
        RECT 5.320 0.695 6.315 0.710 ;
        RECT 5.335 0.675 6.315 0.695 ;
        RECT 5.345 0.655 6.315 0.675 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.195 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.390 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END VPWR
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 7.595 1.585 7.765 2.415 ;
        RECT 8.405 1.585 8.685 2.415 ;
        RECT 7.595 1.415 8.685 1.585 ;
        RECT 8.405 0.905 8.685 1.415 ;
        RECT 7.595 0.735 8.685 0.905 ;
        RECT 7.595 0.315 7.845 0.735 ;
        RECT 8.405 0.315 8.685 0.735 ;
    END
  END COUT
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.335 0.845 2.415 ;
        RECT 1.355 1.565 1.685 2.415 ;
        RECT 1.355 1.335 1.550 1.565 ;
        RECT 0.515 1.065 1.550 1.335 ;
        RECT 0.515 0.315 0.845 1.065 ;
        RECT 1.355 0.825 1.550 1.065 ;
        RECT 1.355 0.315 1.685 0.825 ;
    END
  END SUM
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.135 1.495 0.345 2.635 ;
        RECT 1.015 1.515 1.185 2.635 ;
        RECT 1.855 1.495 2.365 2.635 ;
        RECT 2.770 1.935 2.940 2.355 ;
        RECT 3.190 2.105 3.360 2.635 ;
        RECT 3.530 2.205 4.330 2.375 ;
        RECT 5.240 2.205 5.570 2.635 ;
        RECT 3.530 1.935 3.700 2.205 ;
        RECT 5.835 2.025 6.005 2.355 ;
        RECT 6.175 2.205 6.505 2.635 ;
        RECT 6.675 2.025 6.845 2.355 ;
        RECT 7.055 2.205 7.385 2.635 ;
        RECT 2.580 1.765 3.700 1.935 ;
        RECT 3.870 1.855 7.395 2.025 ;
        RECT 2.580 1.245 2.750 1.765 ;
        RECT 3.870 1.595 4.040 1.855 ;
        RECT 1.720 1.075 2.750 1.245 ;
        RECT 0.135 0.085 0.345 0.885 ;
        RECT 1.015 0.085 1.185 0.885 ;
        RECT 1.855 0.085 2.095 0.885 ;
        RECT 2.580 0.815 2.750 1.075 ;
        RECT 2.920 1.425 4.040 1.595 ;
        RECT 2.920 0.995 3.090 1.425 ;
        RECT 7.225 1.245 7.395 1.855 ;
        RECT 7.935 1.755 8.225 2.635 ;
        RECT 8.855 1.495 9.065 2.635 ;
        RECT 7.225 1.075 8.225 1.245 ;
        RECT 7.225 0.815 7.395 1.075 ;
        RECT 2.580 0.645 3.045 0.815 ;
        RECT 3.215 0.645 5.115 0.815 ;
        RECT 3.215 0.475 3.385 0.645 ;
        RECT 2.270 0.305 3.385 0.475 ;
        RECT 3.555 0.085 3.910 0.465 ;
        RECT 4.080 0.345 4.250 0.645 ;
        RECT 4.920 0.585 5.115 0.645 ;
        RECT 6.705 0.645 7.395 0.815 ;
        RECT 4.420 0.085 4.750 0.465 ;
        RECT 4.920 0.255 5.190 0.585 ;
        RECT 6.705 0.465 6.875 0.645 ;
        RECT 5.385 0.085 5.715 0.465 ;
        RECT 6.175 0.295 6.875 0.465 ;
        RECT 7.055 0.085 7.385 0.465 ;
        RECT 8.015 0.085 8.225 0.565 ;
        RECT 8.855 0.085 9.065 0.885 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
  END
END sky130_fd_sc_hd__ha_4

#--------EOF---------

MACRO sky130_fd_sc_hd__inv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.320 1.075 0.650 1.315 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.210 0.105 1.140 1.015 ;
        RECT 0.210 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 0.720 1.485 1.050 2.465 ;
        RECT 0.820 0.885 1.050 1.485 ;
        RECT 0.720 0.255 1.050 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.340 1.495 0.550 2.635 ;
        RECT 0.320 0.085 0.550 0.905 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
END sky130_fd_sc_hd__inv_1

#--------EOF---------

MACRO sky130_fd_sc_hd__inv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.435 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.105 1.365 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.525 1.485 0.855 2.465 ;
        RECT 0.605 0.885 0.855 1.485 ;
        RECT 0.525 0.255 0.855 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.125 1.495 0.355 2.635 ;
        RECT 1.025 1.495 1.235 2.635 ;
        RECT 0.125 0.085 0.355 0.905 ;
        RECT 1.025 0.085 1.235 0.905 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
END sky130_fd_sc_hd__inv_2

#--------EOF---------

MACRO sky130_fd_sc_hd__inv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 1.735 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.055 0.105 2.245 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.565 1.665 0.895 2.465 ;
        RECT 1.405 1.685 1.735 2.465 ;
        RECT 1.405 1.665 2.170 1.685 ;
        RECT 0.565 1.495 2.170 1.665 ;
        RECT 1.905 0.905 2.170 1.495 ;
        RECT 0.565 0.725 2.170 0.905 ;
        RECT 0.565 0.255 0.895 0.725 ;
        RECT 1.405 0.255 1.735 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.130 1.495 0.395 2.635 ;
        RECT 1.065 1.835 1.235 2.635 ;
        RECT 1.905 2.175 2.115 2.635 ;
        RECT 0.130 0.085 0.395 0.545 ;
        RECT 1.065 0.085 1.235 0.545 ;
        RECT 1.905 0.085 2.155 0.550 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__inv_4

#--------EOF---------

MACRO sky130_fd_sc_hd__inv_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.485000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 2.615 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.055 0.105 3.215 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER li1 ;
        RECT 0.685 1.665 1.015 2.465 ;
        RECT 1.525 1.665 1.855 2.465 ;
        RECT 2.365 1.685 2.695 2.465 ;
        RECT 2.365 1.665 3.135 1.685 ;
        RECT 0.685 1.495 3.135 1.665 ;
        RECT 2.785 0.905 3.135 1.495 ;
        RECT 0.765 0.725 3.135 0.905 ;
        RECT 0.765 0.255 0.935 0.725 ;
        RECT 1.605 0.255 1.775 0.725 ;
        RECT 2.445 0.255 2.615 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.130 1.495 0.425 2.635 ;
        RECT 1.185 1.835 1.355 2.635 ;
        RECT 2.025 1.835 2.195 2.635 ;
        RECT 2.865 2.175 3.035 2.635 ;
        RECT 0.130 0.085 0.395 0.545 ;
        RECT 1.185 0.085 1.355 0.545 ;
        RECT 2.025 0.085 2.195 0.545 ;
        RECT 2.785 0.085 3.035 0.550 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__inv_6

#--------EOF---------

MACRO sky130_fd_sc_hd__inv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 0.680 1.075 3.535 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.170 0.105 4.040 1.015 ;
        RECT 0.170 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 0.680 1.665 1.010 2.465 ;
        RECT 1.520 1.665 1.850 2.465 ;
        RECT 2.360 1.665 2.690 2.465 ;
        RECT 3.200 1.665 3.530 2.465 ;
        RECT 0.085 1.495 4.055 1.665 ;
        RECT 0.085 0.905 0.430 1.495 ;
        RECT 3.735 0.905 4.055 1.495 ;
        RECT 0.085 0.715 4.055 0.905 ;
        RECT 0.680 0.255 1.010 0.715 ;
        RECT 1.520 0.255 1.850 0.715 ;
        RECT 2.360 0.255 2.690 0.715 ;
        RECT 3.200 0.255 3.530 0.715 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.255 1.835 0.510 2.635 ;
        RECT 1.180 1.835 1.350 2.635 ;
        RECT 2.020 1.835 2.190 2.635 ;
        RECT 2.860 1.835 3.030 2.635 ;
        RECT 3.700 1.835 4.000 2.635 ;
        RECT 0.255 0.085 0.510 0.545 ;
        RECT 1.180 0.085 1.350 0.545 ;
        RECT 2.020 0.085 2.190 0.545 ;
        RECT 2.860 0.085 3.030 0.545 ;
        RECT 3.700 0.085 4.005 0.545 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__inv_8

#--------EOF---------

MACRO sky130_fd_sc_hd__inv_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.970000 ;
    PORT
      LAYER li1 ;
        RECT 0.680 1.075 5.270 1.325 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.170 0.105 5.975 1.015 ;
        RECT 0.170 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER li1 ;
        RECT 0.680 1.665 1.010 2.465 ;
        RECT 1.520 1.665 1.850 2.465 ;
        RECT 2.360 1.665 2.690 2.465 ;
        RECT 3.200 1.665 3.530 2.465 ;
        RECT 4.040 1.665 4.370 2.465 ;
        RECT 4.880 1.665 5.210 2.465 ;
        RECT 0.085 1.495 5.895 1.665 ;
        RECT 0.085 0.905 0.510 1.495 ;
        RECT 5.545 0.905 5.895 1.495 ;
        RECT 0.085 0.715 5.895 0.905 ;
        RECT 0.680 0.255 1.010 0.715 ;
        RECT 1.520 0.255 1.850 0.715 ;
        RECT 2.360 0.255 2.690 0.715 ;
        RECT 3.200 0.255 3.530 0.715 ;
        RECT 4.040 0.255 4.370 0.715 ;
        RECT 4.880 0.255 5.210 0.715 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.255 1.835 0.510 2.635 ;
        RECT 1.180 1.835 1.350 2.635 ;
        RECT 2.020 1.835 2.190 2.635 ;
        RECT 2.860 1.835 3.030 2.635 ;
        RECT 3.700 1.835 3.870 2.635 ;
        RECT 4.540 1.835 4.710 2.635 ;
        RECT 5.555 1.835 5.895 2.635 ;
        RECT 0.255 0.085 0.510 0.545 ;
        RECT 1.180 0.085 1.350 0.545 ;
        RECT 2.020 0.085 2.190 0.545 ;
        RECT 2.860 0.085 3.030 0.545 ;
        RECT 3.700 0.085 3.870 0.545 ;
        RECT 4.540 0.085 4.710 0.545 ;
        RECT 5.555 0.085 5.895 0.545 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
END sky130_fd_sc_hd__inv_12

#--------EOF---------

MACRO sky130_fd_sc_hd__inv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__inv_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.960000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 5.525 1.315 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.070 0.105 7.300 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER li1 ;
        RECT 0.580 1.665 0.910 2.465 ;
        RECT 1.420 1.665 1.750 2.465 ;
        RECT 2.260 1.665 2.590 2.465 ;
        RECT 3.100 1.665 3.430 2.465 ;
        RECT 3.940 1.665 4.270 2.465 ;
        RECT 4.780 1.665 5.110 2.465 ;
        RECT 5.620 1.665 5.950 2.465 ;
        RECT 6.460 1.665 6.790 2.465 ;
        RECT 0.580 1.495 6.790 1.665 ;
        RECT 6.460 0.905 6.790 1.495 ;
        RECT 0.580 0.715 6.790 0.905 ;
        RECT 0.580 0.255 0.910 0.715 ;
        RECT 1.420 0.255 1.750 0.715 ;
        RECT 2.260 0.255 2.590 0.715 ;
        RECT 3.100 0.255 3.430 0.715 ;
        RECT 3.940 0.255 4.270 0.715 ;
        RECT 4.780 0.255 5.110 0.715 ;
        RECT 5.620 0.255 5.950 0.715 ;
        RECT 6.460 0.255 6.790 0.715 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.200 1.485 0.410 2.635 ;
        RECT 1.080 1.835 1.250 2.635 ;
        RECT 1.920 1.835 2.090 2.635 ;
        RECT 2.760 1.835 2.930 2.635 ;
        RECT 3.600 1.835 3.770 2.635 ;
        RECT 4.440 1.835 4.610 2.635 ;
        RECT 5.280 1.835 5.450 2.635 ;
        RECT 6.120 1.835 6.290 2.635 ;
        RECT 6.960 1.835 7.170 2.635 ;
        RECT 0.180 0.085 0.410 0.885 ;
        RECT 1.080 0.085 1.250 0.545 ;
        RECT 1.920 0.085 2.090 0.545 ;
        RECT 2.760 0.085 2.930 0.545 ;
        RECT 3.600 0.085 3.770 0.545 ;
        RECT 4.440 0.085 4.610 0.545 ;
        RECT 5.280 0.085 5.450 0.545 ;
        RECT 6.120 0.085 6.290 0.545 ;
        RECT 6.960 0.085 7.170 0.885 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
END sky130_fd_sc_hd__inv_16

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_bleeder_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_bleeder_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN SHORT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.270000 ;
    PORT
      LAYER li1 ;
        RECT 0.275 1.040 1.975 1.730 ;
    END
  END SHORT
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.195 0.395 2.565 1.015 ;
        RECT 0.195 0.085 0.315 0.395 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.285 0.085 0.615 0.870 ;
        RECT 2.145 0.540 2.475 2.635 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_bleeder_1

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.985 1.275 1.355 ;
    END
  END A
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 1.310 2.340 ;
        RECT 0.550 2.080 0.840 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.375 0.885 ;
        RECT 1.065 -0.085 1.235 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.560 0.355 2.465 ;
        RECT 0.085 0.760 0.255 1.560 ;
        RECT 0.085 0.255 0.345 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.525 1.875 0.855 2.465 ;
        RECT 1.035 1.705 1.205 2.465 ;
        RECT 0.540 1.535 1.205 1.705 ;
        RECT 0.540 1.390 0.710 1.535 ;
        RECT 0.425 1.060 0.710 1.390 ;
        RECT 0.540 0.805 0.710 1.060 ;
        RECT 0.540 0.635 1.205 0.805 ;
        RECT 0.525 0.085 0.855 0.465 ;
        RECT 1.035 0.255 1.205 0.635 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.610 2.125 0.780 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_1

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.745 0.785 1.240 ;
    END
  END A
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 1.770 2.340 ;
        RECT 0.550 2.080 0.840 2.140 ;
        RECT 1.435 2.080 1.725 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.835 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER li1 ;
        RECT 1.060 1.970 1.245 2.435 ;
        RECT 1.060 1.750 1.725 1.970 ;
        RECT 1.385 0.825 1.725 1.750 ;
        RECT 1.040 0.655 1.725 0.825 ;
        RECT 1.040 0.255 1.245 0.655 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.085 1.580 0.355 2.435 ;
        RECT 0.525 1.855 0.855 2.465 ;
        RECT 1.415 2.140 1.750 2.465 ;
        RECT 0.085 1.410 1.215 1.580 ;
        RECT 0.085 0.585 0.255 1.410 ;
        RECT 0.965 0.995 1.215 1.410 ;
        RECT 0.085 0.255 0.345 0.585 ;
        RECT 0.555 0.085 0.830 0.565 ;
        RECT 1.415 0.085 1.750 0.485 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.610 2.125 0.780 2.295 ;
        RECT 1.495 2.140 1.665 2.310 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_2

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.755 0.775 1.325 ;
    END
  END A
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 2.690 2.340 ;
        RECT 0.550 2.080 0.840 2.140 ;
        RECT 1.435 2.080 1.725 2.140 ;
        RECT 2.315 2.080 2.605 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.745 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER li1 ;
        RECT 1.025 2.005 1.265 2.465 ;
        RECT 1.025 2.000 1.325 2.005 ;
        RECT 1.025 1.980 1.330 2.000 ;
        RECT 1.025 1.975 1.370 1.980 ;
        RECT 1.025 1.970 1.385 1.975 ;
        RECT 1.025 1.965 1.390 1.970 ;
        RECT 1.935 1.965 2.165 2.465 ;
        RECT 1.025 1.835 2.165 1.965 ;
        RECT 1.185 1.825 2.165 1.835 ;
        RECT 1.195 1.820 2.165 1.825 ;
        RECT 1.205 1.815 2.165 1.820 ;
        RECT 1.215 1.805 2.165 1.815 ;
        RECT 1.245 1.785 2.165 1.805 ;
        RECT 1.270 1.750 2.165 1.785 ;
        RECT 1.905 1.585 2.165 1.750 ;
        RECT 1.905 1.415 2.660 1.585 ;
        RECT 2.255 0.905 2.660 1.415 ;
        RECT 1.010 0.735 2.660 0.905 ;
        RECT 1.010 0.345 1.305 0.735 ;
        RECT 1.905 0.345 2.165 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.085 1.665 0.355 2.465 ;
        RECT 0.525 1.835 0.855 2.465 ;
        RECT 1.435 2.140 1.765 2.465 ;
        RECT 2.335 1.765 2.620 2.465 ;
        RECT 0.085 1.495 1.115 1.665 ;
        RECT 0.085 0.585 0.255 1.495 ;
        RECT 0.945 1.245 1.115 1.495 ;
        RECT 0.945 1.075 2.085 1.245 ;
        RECT 0.085 0.255 0.385 0.585 ;
        RECT 0.555 0.085 0.830 0.565 ;
        RECT 1.475 0.085 1.730 0.565 ;
        RECT 2.335 0.085 2.615 0.565 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.610 2.125 0.780 2.295 ;
        RECT 1.495 2.140 1.665 2.310 ;
        RECT 2.375 2.125 2.545 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_4

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.715 0.400 1.325 ;
    END
  END A
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 4.990 2.340 ;
        RECT 0.115 2.080 0.405 2.140 ;
        RECT 0.975 2.080 1.265 2.140 ;
        RECT 1.830 2.080 2.120 2.140 ;
        RECT 2.680 2.080 2.970 2.140 ;
        RECT 3.560 2.080 3.850 2.140 ;
        RECT 4.420 2.080 4.710 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.820 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER li1 ;
        RECT 1.420 1.735 1.680 2.460 ;
        RECT 2.280 1.735 2.540 2.460 ;
        RECT 3.140 1.735 3.400 2.460 ;
        RECT 4.000 1.735 4.260 2.460 ;
        RECT 1.420 1.495 4.730 1.735 ;
        RECT 3.760 0.905 4.730 1.495 ;
        RECT 1.420 0.735 4.730 0.905 ;
        RECT 1.420 0.280 1.680 0.735 ;
        RECT 2.280 0.280 2.540 0.735 ;
        RECT 3.140 0.280 3.400 0.735 ;
        RECT 4.000 0.280 4.260 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.095 1.525 0.390 2.465 ;
        RECT 0.570 1.325 0.820 2.460 ;
        RECT 0.990 1.525 1.250 2.465 ;
        RECT 1.850 1.905 2.110 2.465 ;
        RECT 2.710 1.905 2.970 2.465 ;
        RECT 3.570 1.905 3.830 2.465 ;
        RECT 4.430 1.905 4.725 2.465 ;
        RECT 0.570 1.075 3.590 1.325 ;
        RECT 0.145 0.085 0.390 0.545 ;
        RECT 0.570 0.265 0.820 1.075 ;
        RECT 0.990 0.085 1.250 0.610 ;
        RECT 1.850 0.085 2.110 0.565 ;
        RECT 2.710 0.085 2.970 0.565 ;
        RECT 3.570 0.085 3.830 0.565 ;
        RECT 4.430 0.085 4.730 0.565 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.175 2.125 0.345 2.295 ;
        RECT 1.035 2.125 1.205 2.295 ;
        RECT 1.890 2.125 2.060 2.295 ;
        RECT 2.740 2.125 2.910 2.295 ;
        RECT 3.620 2.125 3.790 2.295 ;
        RECT 4.480 2.125 4.650 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_8

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_clkbufkapwr_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkbufkapwr_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.400 1.325 ;
    END
  END A
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 9.130 2.340 ;
        RECT 0.115 2.080 0.405 2.140 ;
        RECT 0.975 2.080 1.265 2.140 ;
        RECT 1.830 2.080 2.120 2.140 ;
        RECT 2.680 2.080 2.970 2.140 ;
        RECT 3.560 2.080 3.850 2.140 ;
        RECT 4.420 2.080 4.710 2.140 ;
        RECT 5.275 2.080 5.565 2.140 ;
        RECT 6.135 2.080 6.425 2.140 ;
        RECT 6.990 2.080 7.280 2.140 ;
        RECT 7.840 2.080 8.130 2.140 ;
        RECT 8.720 2.080 9.010 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.110 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.390 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER li1 ;
        RECT 2.315 1.735 2.540 2.460 ;
        RECT 3.140 1.735 3.400 2.460 ;
        RECT 4.000 1.735 4.260 2.460 ;
        RECT 4.860 1.735 5.120 2.460 ;
        RECT 5.705 1.735 5.965 2.460 ;
        RECT 6.565 1.735 6.825 2.460 ;
        RECT 7.425 1.735 7.685 2.460 ;
        RECT 2.315 1.720 7.685 1.735 ;
        RECT 8.295 1.720 8.585 2.460 ;
        RECT 2.315 1.495 9.025 1.720 ;
        RECT 7.860 0.905 9.025 1.495 ;
        RECT 2.280 0.735 9.025 0.905 ;
        RECT 2.280 0.280 2.540 0.735 ;
        RECT 3.140 0.280 3.400 0.735 ;
        RECT 4.000 0.280 4.260 0.735 ;
        RECT 4.845 0.280 5.120 0.735 ;
        RECT 5.705 0.280 5.965 0.735 ;
        RECT 6.565 0.280 6.825 0.735 ;
        RECT 7.425 0.280 7.685 0.735 ;
        RECT 8.295 0.280 8.555 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.095 1.495 0.425 2.465 ;
        RECT 0.595 1.325 0.785 2.465 ;
        RECT 0.955 1.495 1.285 2.465 ;
        RECT 1.455 1.325 1.645 2.460 ;
        RECT 1.815 1.495 2.145 2.465 ;
        RECT 2.710 1.905 2.970 2.465 ;
        RECT 3.570 1.905 3.830 2.465 ;
        RECT 4.430 1.905 4.690 2.465 ;
        RECT 5.290 1.905 5.535 2.465 ;
        RECT 6.150 1.905 6.395 2.465 ;
        RECT 7.010 1.905 7.255 2.465 ;
        RECT 7.870 1.905 8.125 2.465 ;
        RECT 8.755 1.890 9.025 2.465 ;
        RECT 0.595 1.075 7.690 1.325 ;
        RECT 0.085 0.085 0.390 0.595 ;
        RECT 0.595 0.265 0.820 1.075 ;
        RECT 0.990 0.085 1.250 0.610 ;
        RECT 1.430 0.265 1.680 1.075 ;
        RECT 1.850 0.085 2.110 0.645 ;
        RECT 2.710 0.085 2.970 0.565 ;
        RECT 3.570 0.085 3.830 0.565 ;
        RECT 4.430 0.085 4.675 0.565 ;
        RECT 5.290 0.085 5.535 0.565 ;
        RECT 6.145 0.085 6.395 0.565 ;
        RECT 7.005 0.085 7.255 0.565 ;
        RECT 7.865 0.085 8.125 0.565 ;
        RECT 8.725 0.085 9.025 0.565 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 0.175 2.125 0.345 2.295 ;
        RECT 1.035 2.125 1.205 2.295 ;
        RECT 1.890 2.125 2.060 2.295 ;
        RECT 2.740 2.125 2.910 2.295 ;
        RECT 3.620 2.125 3.790 2.295 ;
        RECT 4.480 2.125 4.650 2.295 ;
        RECT 5.335 2.125 5.505 2.295 ;
        RECT 6.195 2.125 6.365 2.295 ;
        RECT 7.050 2.125 7.220 2.295 ;
        RECT 7.900 2.125 8.070 2.295 ;
        RECT 8.780 2.125 8.950 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_clkbufkapwr_16

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.315000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.375 0.325 1.325 ;
    END
  END A
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 1.310 2.340 ;
        RECT 0.095 2.080 0.385 2.140 ;
        RECT 0.995 2.080 1.285 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.336000 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.290 0.765 2.465 ;
        RECT 0.595 0.945 1.295 1.290 ;
        RECT 0.590 0.760 1.295 0.945 ;
        RECT 0.590 0.255 0.840 0.760 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 0.420 0.105 1.375 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.085 1.665 0.425 2.465 ;
        RECT 0.935 1.665 1.295 2.465 ;
        RECT 1.010 0.085 1.295 0.590 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.155 2.125 0.325 2.295 ;
        RECT 1.055 2.125 1.225 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_1

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.576000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.065 1.305 1.290 ;
    END
  END A
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 1.770 2.340 ;
        RECT 0.540 2.080 0.830 2.140 ;
        RECT 1.440 2.080 1.730 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.662600 ;
    PORT
      LAYER li1 ;
        RECT 0.155 1.630 0.375 2.435 ;
        RECT 1.045 1.630 1.235 2.435 ;
        RECT 0.155 1.460 1.755 1.630 ;
        RECT 1.475 0.895 1.755 1.460 ;
        RECT 1.025 0.725 1.755 0.895 ;
        RECT 1.025 0.280 1.250 0.725 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 0.470 0.105 1.835 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.545 1.800 0.875 2.465 ;
        RECT 1.405 1.800 1.735 2.465 ;
        RECT 0.560 0.085 0.855 0.610 ;
        RECT 1.420 0.085 1.750 0.555 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.600 2.125 0.770 2.295 ;
        RECT 1.500 2.125 1.670 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_2

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.152000 ;
    PORT
      LAYER li1 ;
        RECT 0.445 1.065 2.660 1.290 ;
    END
  END A
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 3.150 2.340 ;
        RECT 0.135 2.080 0.425 2.140 ;
        RECT 0.995 2.080 1.285 2.140 ;
        RECT 1.895 2.080 2.185 2.140 ;
        RECT 2.775 2.080 3.065 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.075200 ;
    PORT
      LAYER li1 ;
        RECT 0.645 1.630 0.815 2.435 ;
        RECT 1.505 1.630 1.675 2.435 ;
        RECT 2.365 1.630 2.535 2.435 ;
        RECT 0.105 1.460 3.135 1.630 ;
        RECT 0.105 0.895 0.275 1.460 ;
        RECT 2.835 0.895 3.135 1.460 ;
        RECT 0.105 0.725 3.135 0.895 ;
        RECT 1.030 0.280 1.290 0.725 ;
        RECT 1.890 0.280 2.145 0.725 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 0.410 0.105 2.835 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.135 1.800 0.465 2.465 ;
        RECT 0.995 1.800 1.325 2.465 ;
        RECT 1.855 1.800 2.185 2.465 ;
        RECT 2.715 1.800 3.045 2.465 ;
        RECT 0.565 0.085 0.860 0.555 ;
        RECT 1.460 0.085 1.720 0.555 ;
        RECT 2.315 0.085 2.615 0.555 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.195 2.125 0.365 2.295 ;
        RECT 1.055 2.125 1.225 2.295 ;
        RECT 1.955 2.125 2.125 2.295 ;
        RECT 2.835 2.125 3.005 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_4

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.304000 ;
    PORT
      LAYER li1 ;
        RECT 0.455 1.035 4.865 1.290 ;
    END
  END A
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 5.910 2.340 ;
        RECT 0.070 2.080 0.360 2.140 ;
        RECT 0.930 2.080 1.220 2.140 ;
        RECT 1.830 2.080 2.120 2.140 ;
        RECT 2.710 2.080 3.000 2.140 ;
        RECT 3.435 2.080 3.725 2.140 ;
        RECT 4.295 2.080 4.585 2.140 ;
        RECT 5.195 2.080 5.485 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150 -0.085 0.320 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.090400 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.630 0.765 2.435 ;
        RECT 1.440 1.630 1.610 2.435 ;
        RECT 2.280 1.630 2.450 2.435 ;
        RECT 3.120 1.630 3.290 2.435 ;
        RECT 3.960 1.630 4.130 2.435 ;
        RECT 4.800 1.630 4.970 2.435 ;
        RECT 0.115 1.460 5.440 1.630 ;
        RECT 0.115 0.865 0.285 1.460 ;
        RECT 5.170 0.865 5.440 1.460 ;
        RECT 0.115 0.695 5.440 0.865 ;
        RECT 1.535 0.280 1.725 0.695 ;
        RECT 2.395 0.280 2.585 0.695 ;
        RECT 3.255 0.280 3.445 0.695 ;
        RECT 4.115 0.280 4.305 0.695 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 0.945 0.105 4.895 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.095 1.800 0.425 2.465 ;
        RECT 0.940 1.800 1.270 2.465 ;
        RECT 1.780 1.800 2.110 2.465 ;
        RECT 2.620 1.800 2.950 2.465 ;
        RECT 3.460 1.800 3.790 2.465 ;
        RECT 4.300 1.800 4.630 2.465 ;
        RECT 5.140 1.800 5.470 2.465 ;
        RECT 1.035 0.085 1.365 0.525 ;
        RECT 1.895 0.085 2.225 0.525 ;
        RECT 2.755 0.085 3.085 0.525 ;
        RECT 3.615 0.085 3.945 0.525 ;
        RECT 4.475 0.085 4.805 0.525 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.130 2.125 0.300 2.295 ;
        RECT 0.990 2.125 1.160 2.295 ;
        RECT 1.890 2.125 2.060 2.295 ;
        RECT 2.770 2.125 2.940 2.295 ;
        RECT 3.495 2.125 3.665 2.295 ;
        RECT 4.355 2.125 4.525 2.295 ;
        RECT 5.255 2.125 5.425 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_8

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.608000 ;
    PORT
      LAYER met1 ;
        RECT 1.465 1.260 2.215 1.305 ;
        RECT 9.285 1.260 10.035 1.305 ;
        RECT 1.465 1.120 10.035 1.260 ;
        RECT 1.465 1.075 2.215 1.120 ;
        RECT 9.285 1.075 10.035 1.120 ;
    END
  END A
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 10.970 2.340 ;
        RECT 0.070 2.080 0.360 2.140 ;
        RECT 0.930 2.080 1.220 2.140 ;
        RECT 1.830 2.080 2.120 2.140 ;
        RECT 2.710 2.080 3.000 2.140 ;
        RECT 3.630 2.080 3.920 2.140 ;
        RECT 4.490 2.080 4.780 2.140 ;
        RECT 5.390 2.080 5.680 2.140 ;
        RECT 6.310 2.080 6.600 2.140 ;
        RECT 7.170 2.080 7.460 2.140 ;
        RECT 8.070 2.080 8.360 2.140 ;
        RECT 8.900 2.080 9.190 2.140 ;
        RECT 9.760 2.080 10.050 2.140 ;
        RECT 10.660 2.080 10.950 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.520900 ;
    PORT
      LAYER li1 ;
        RECT 0.615 1.665 0.785 2.465 ;
        RECT 1.475 1.665 1.645 2.465 ;
        RECT 2.335 1.665 2.505 2.465 ;
        RECT 3.195 1.665 3.365 2.465 ;
        RECT 4.055 1.665 4.225 2.465 ;
        RECT 5.080 1.665 5.250 2.465 ;
        RECT 5.965 1.665 6.135 2.465 ;
        RECT 6.825 1.665 6.995 2.465 ;
        RECT 7.685 1.665 7.855 2.465 ;
        RECT 8.545 1.665 8.715 2.465 ;
        RECT 9.405 1.665 9.575 2.465 ;
        RECT 10.265 1.665 10.435 2.465 ;
        RECT 0.615 1.455 10.480 1.665 ;
        RECT 2.325 1.415 8.755 1.455 ;
        RECT 2.325 0.280 2.550 1.415 ;
        RECT 3.155 0.280 3.410 1.415 ;
        RECT 4.015 0.280 4.255 1.415 ;
        RECT 4.905 0.280 5.255 1.415 ;
        RECT 5.925 0.280 6.175 1.415 ;
        RECT 6.785 0.280 7.035 1.415 ;
        RECT 7.645 0.280 7.895 1.415 ;
        RECT 8.505 0.280 8.755 1.415 ;
    END
  END Y
  OBS
      LAYER pwell ;
        RECT 1.735 0.105 9.315 0.785 ;
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.110 1.495 0.440 2.465 ;
        RECT 0.965 1.835 1.295 2.465 ;
        RECT 1.825 1.835 2.155 2.465 ;
        RECT 2.685 1.835 3.015 2.465 ;
        RECT 3.545 1.835 3.875 2.465 ;
        RECT 4.425 1.835 4.755 2.465 ;
        RECT 5.450 1.835 5.780 2.465 ;
        RECT 6.315 1.835 6.645 2.465 ;
        RECT 7.175 1.835 7.505 2.465 ;
        RECT 8.035 1.835 8.365 2.465 ;
        RECT 8.895 1.835 9.225 2.465 ;
        RECT 9.755 1.835 10.085 2.465 ;
        RECT 10.610 1.835 10.940 2.465 ;
        RECT 0.345 0.895 2.155 1.275 ;
        RECT 8.930 0.895 10.710 1.275 ;
        RECT 1.855 0.085 2.125 0.610 ;
        RECT 2.720 0.085 2.985 0.610 ;
        RECT 3.580 0.085 3.845 0.610 ;
        RECT 4.465 0.085 4.730 0.610 ;
        RECT 5.490 0.085 5.755 0.610 ;
        RECT 6.350 0.085 6.575 0.610 ;
        RECT 7.210 0.085 7.475 0.610 ;
        RECT 8.070 0.085 8.335 0.610 ;
        RECT 8.930 0.085 9.195 0.610 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 0.130 2.125 0.300 2.295 ;
        RECT 0.990 2.125 1.160 2.295 ;
        RECT 1.890 2.125 2.060 2.295 ;
        RECT 2.770 2.125 2.940 2.295 ;
        RECT 3.690 2.125 3.860 2.295 ;
        RECT 4.550 2.125 4.720 2.295 ;
        RECT 5.450 2.125 5.620 2.295 ;
        RECT 6.370 2.125 6.540 2.295 ;
        RECT 7.230 2.125 7.400 2.295 ;
        RECT 8.130 2.125 8.300 2.295 ;
        RECT 8.960 2.125 9.130 2.295 ;
        RECT 9.820 2.125 9.990 2.295 ;
        RECT 10.720 2.125 10.890 2.295 ;
        RECT 1.525 1.105 1.695 1.275 ;
        RECT 1.985 1.105 2.155 1.275 ;
        RECT 9.345 1.105 9.515 1.275 ;
        RECT 9.805 1.105 9.975 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_clkinvkapwr_16

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_decapkapwr_3
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 1.310 2.340 ;
        RECT 0.085 2.080 1.295 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.375 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.085 1.545 1.295 2.465 ;
        RECT 0.085 0.835 0.605 1.375 ;
        RECT 0.775 1.005 1.295 1.545 ;
        RECT 0.085 0.085 1.295 0.835 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 2.125 0.315 2.295 ;
        RECT 0.605 2.125 0.775 2.295 ;
        RECT 1.065 2.125 1.235 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_3

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_decapkapwr_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 1.770 2.340 ;
        RECT 0.085 2.080 1.755 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.835 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.085 1.545 1.755 2.465 ;
        RECT 0.085 0.855 0.835 1.375 ;
        RECT 1.005 1.025 1.755 1.545 ;
        RECT 0.085 0.085 1.755 0.855 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 2.125 0.315 2.295 ;
        RECT 0.605 2.125 0.775 2.295 ;
        RECT 1.065 2.125 1.235 2.295 ;
        RECT 1.525 2.125 1.695 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_4

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_decapkapwr_6
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 2.690 2.340 ;
        RECT 0.085 2.080 2.675 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.755 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.085 1.545 2.675 2.465 ;
        RECT 0.085 0.855 1.295 1.375 ;
        RECT 1.465 1.025 2.675 1.545 ;
        RECT 0.085 0.085 2.675 0.855 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 2.125 0.315 2.295 ;
        RECT 0.605 2.125 0.775 2.295 ;
        RECT 1.065 2.125 1.235 2.295 ;
        RECT 1.525 2.125 1.695 2.295 ;
        RECT 1.985 2.125 2.155 2.295 ;
        RECT 2.445 2.125 2.615 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_6

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_decapkapwr_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 3.610 2.340 ;
        RECT 0.085 2.080 3.595 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.675 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.545 3.595 2.465 ;
        RECT 0.085 0.855 1.735 1.375 ;
        RECT 1.905 1.025 3.595 1.545 ;
        RECT 0.085 0.085 3.595 0.855 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 2.125 0.315 2.295 ;
        RECT 0.605 2.125 0.775 2.295 ;
        RECT 1.065 2.125 1.235 2.295 ;
        RECT 1.525 2.125 1.695 2.295 ;
        RECT 1.985 2.125 2.155 2.295 ;
        RECT 2.445 2.125 2.615 2.295 ;
        RECT 2.905 2.125 3.075 2.295 ;
        RECT 3.365 2.125 3.535 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_8

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_decapkapwr_12
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_decapkapwr_12 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 5.450 2.340 ;
        RECT 0.085 2.080 5.435 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.515 0.915 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.085 1.545 5.430 2.465 ;
        RECT 0.085 0.855 2.665 1.375 ;
        RECT 2.835 1.025 5.430 1.545 ;
        RECT 0.085 0.085 5.430 0.855 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 2.125 0.315 2.295 ;
        RECT 0.605 2.125 0.775 2.295 ;
        RECT 1.065 2.125 1.235 2.295 ;
        RECT 1.525 2.125 1.695 2.295 ;
        RECT 1.985 2.125 2.155 2.295 ;
        RECT 2.445 2.125 2.615 2.295 ;
        RECT 2.905 2.125 3.075 2.295 ;
        RECT 3.365 2.125 3.535 2.295 ;
        RECT 3.825 2.125 3.995 2.295 ;
        RECT 4.285 2.125 4.455 2.295 ;
        RECT 4.745 2.125 4.915 2.295 ;
        RECT 5.205 2.125 5.375 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_decapkapwr_12

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_inputiso0n_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso0n_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.325 0.365 1.685 ;
        RECT 0.100 1.075 0.775 1.325 ;
    END
  END A
  PIN SLEEP_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.075 1.335 1.325 ;
    END
  END SLEEP_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.145 0.925 2.095 1.015 ;
        RECT 0.165 0.105 2.095 0.925 ;
        RECT 0.165 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.657000 ;
    PORT
      LAYER li1 ;
        RECT 1.755 1.915 2.215 2.465 ;
        RECT 1.965 0.545 2.215 1.915 ;
        RECT 1.655 0.255 2.215 0.545 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.285 1.965 0.565 2.635 ;
        RECT 0.735 1.745 1.035 2.295 ;
        RECT 1.235 1.915 1.565 2.635 ;
        RECT 0.735 1.575 1.675 1.745 ;
        RECT 1.505 1.325 1.675 1.575 ;
        RECT 1.505 0.995 1.795 1.325 ;
        RECT 1.505 0.905 1.675 0.995 ;
        RECT 0.285 0.715 1.675 0.905 ;
        RECT 0.285 0.355 0.615 0.715 ;
        RECT 1.235 0.085 1.485 0.545 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso0n_1

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_inputiso0p_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso0p_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.480 1.645 2.175 1.955 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.445 1.615 ;
    END
  END SLEEP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.825 0.785 2.755 1.015 ;
        RECT 0.005 0.105 2.755 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 2.350 1.580 2.655 2.365 ;
        RECT 2.480 0.775 2.655 1.580 ;
        RECT 2.415 0.255 2.655 0.775 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.175 2.015 0.345 2.445 ;
        RECT 0.515 2.185 0.845 2.635 ;
        RECT 0.175 1.785 0.850 2.015 ;
        RECT 0.615 1.135 0.850 1.785 ;
        RECT 1.020 1.475 1.305 2.420 ;
        RECT 1.485 2.165 2.170 2.635 ;
        RECT 1.020 1.325 1.880 1.475 ;
        RECT 1.020 1.305 2.305 1.325 ;
        RECT 0.615 0.805 1.150 1.135 ;
        RECT 1.320 0.945 2.305 1.305 ;
        RECT 0.615 0.655 0.835 0.805 ;
        RECT 0.090 0.085 0.425 0.590 ;
        RECT 0.595 0.280 0.835 0.655 ;
        RECT 1.320 0.610 1.490 0.945 ;
        RECT 1.115 0.415 1.490 0.610 ;
        RECT 1.115 0.270 1.285 0.415 ;
        RECT 1.850 0.085 2.245 0.580 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso0p_1

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_inputiso1n_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso1n_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.540 2.085 1.735 2.415 ;
    END
  END A
  PIN SLEEP_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.425 1.325 ;
    END
  END SLEEP_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.810 0.815 2.755 1.015 ;
        RECT 0.005 0.135 2.755 0.815 ;
        RECT 0.150 -0.085 0.320 0.135 ;
        RECT 1.810 0.105 2.755 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.495 2.675 2.465 ;
        RECT 2.505 0.760 2.675 1.495 ;
        RECT 2.405 0.415 2.675 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 0.595 1.325 0.765 1.885 ;
        RECT 0.990 1.665 1.410 1.915 ;
        RECT 1.915 1.835 2.195 2.635 ;
        RECT 0.990 1.495 2.235 1.665 ;
        RECT 2.065 1.325 2.235 1.495 ;
        RECT 0.595 0.995 1.335 1.325 ;
        RECT 2.065 0.995 2.295 1.325 ;
        RECT 0.595 0.905 0.845 0.995 ;
        RECT 0.110 0.735 0.845 0.905 ;
        RECT 2.065 0.825 2.235 0.995 ;
        RECT 0.110 0.265 0.420 0.735 ;
        RECT 1.495 0.655 2.235 0.825 ;
        RECT 0.590 0.085 1.325 0.565 ;
        RECT 1.495 0.305 1.665 0.655 ;
        RECT 1.835 0.085 2.215 0.485 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso1n_1

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_inputiso1p_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputiso1p_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.500 1.325 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.010 0.765 1.275 1.325 ;
    END
  END SLEEP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.055 0.785 1.985 1.015 ;
        RECT 0.150 0.105 1.985 0.785 ;
        RECT 0.150 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.509000 ;
    PORT
      LAYER li1 ;
        RECT 1.645 1.845 2.180 2.465 ;
        RECT 1.865 0.825 2.180 1.845 ;
        RECT 1.565 0.255 2.180 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.270 1.665 0.660 1.840 ;
        RECT 1.145 1.835 1.475 2.635 ;
        RECT 0.270 1.495 1.695 1.665 ;
        RECT 0.670 0.595 0.840 1.495 ;
        RECT 1.525 0.995 1.695 1.495 ;
        RECT 0.250 0.085 0.490 0.595 ;
        RECT 0.670 0.265 0.950 0.595 ;
        RECT 1.180 0.085 1.395 0.595 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_inputiso1p_1

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_inputisolatch_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_inputisolatch_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.750 0.765 2.125 1.095 ;
    END
  END D
  PIN SLEEP_B
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.145500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.985 0.330 1.625 ;
    END
  END SLEEP_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.725 2.285 0.785 ;
        RECT 3.705 0.725 5.055 1.015 ;
        RECT 0.005 0.105 5.055 0.725 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 4.690 1.670 4.975 2.455 ;
        RECT 4.805 0.745 4.975 1.670 ;
        RECT 4.690 0.415 4.975 0.745 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 1.015 2.085 1.185 2.465 ;
        RECT 1.455 2.255 1.850 2.635 ;
        RECT 2.310 2.255 3.185 2.425 ;
        RECT 1.015 1.965 2.845 2.085 ;
        RECT 0.175 1.795 0.780 1.965 ;
        RECT 0.610 1.460 0.780 1.795 ;
        RECT 0.980 1.915 2.845 1.965 ;
        RECT 0.980 1.825 1.185 1.915 ;
        RECT 0.610 1.130 0.810 1.460 ;
        RECT 0.610 0.805 0.780 1.130 ;
        RECT 0.175 0.635 0.780 0.805 ;
        RECT 0.980 0.910 1.150 1.825 ;
        RECT 1.320 1.525 2.335 1.695 ;
        RECT 1.320 1.240 1.490 1.525 ;
        RECT 2.050 1.355 2.335 1.525 ;
        RECT 2.505 1.575 2.845 1.915 ;
        RECT 2.505 1.035 2.675 1.575 ;
        RECT 3.015 1.325 3.185 2.255 ;
        RECT 3.355 2.135 3.525 2.635 ;
        RECT 3.835 1.865 4.125 2.435 ;
        RECT 3.420 1.535 4.125 1.865 ;
        RECT 4.295 1.570 4.465 2.635 ;
        RECT 3.015 1.165 3.780 1.325 ;
        RECT 0.980 0.740 1.185 0.910 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 0.740 ;
        RECT 2.295 0.705 2.675 1.035 ;
        RECT 2.870 0.995 3.780 1.165 ;
        RECT 2.870 0.535 3.040 0.995 ;
        RECT 3.950 0.745 4.125 1.535 ;
        RECT 1.455 0.085 1.785 0.465 ;
        RECT 2.380 0.365 3.040 0.535 ;
        RECT 3.265 0.085 3.595 0.530 ;
        RECT 3.835 0.415 4.125 0.745 ;
        RECT 4.295 0.085 4.465 0.715 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_inputisolatch_1

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_isobufsrc_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 0.725 0.325 1.325 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.960 1.065 1.325 1.325 ;
    END
  END SLEEP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.725 0.785 2.075 1.015 ;
        RECT 0.240 0.105 2.075 0.785 ;
        RECT 0.240 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.435500 ;
    PORT
      LAYER li1 ;
        RECT 1.655 1.850 2.215 2.465 ;
        RECT 2.035 0.895 2.215 1.850 ;
        RECT 1.235 0.725 2.215 0.895 ;
        RECT 1.235 0.255 1.565 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.415 1.680 0.675 1.905 ;
        RECT 0.875 1.855 1.205 2.635 ;
        RECT 0.415 1.510 1.705 1.680 ;
        RECT 0.495 0.545 0.675 1.510 ;
        RECT 1.535 1.245 1.705 1.510 ;
        RECT 1.535 1.075 1.865 1.245 ;
        RECT 0.330 0.370 0.675 0.545 ;
        RECT 0.855 0.085 1.065 0.895 ;
        RECT 1.735 0.085 2.120 0.555 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_1

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_isobufsrc_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.910 1.275 3.125 1.965 ;
        RECT 2.600 1.065 3.125 1.275 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.480 1.065 0.920 1.275 ;
    END
  END SLEEP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.335 3.155 1.015 ;
        RECT 0.010 0.105 2.215 0.335 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.621000 ;
    PORT
      LAYER li1 ;
        RECT 1.415 0.895 1.665 2.125 ;
        RECT 0.535 0.725 1.705 0.895 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 1.375 0.255 1.705 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.655 0.405 2.465 ;
        RECT 0.575 1.825 0.825 2.635 ;
        RECT 0.995 2.295 2.125 2.465 ;
        RECT 0.995 1.655 1.245 2.295 ;
        RECT 0.085 1.445 1.245 1.655 ;
        RECT 1.835 1.890 2.125 2.295 ;
        RECT 1.835 1.445 2.090 1.890 ;
        RECT 2.395 1.615 2.565 2.460 ;
        RECT 2.775 2.145 3.025 2.635 ;
        RECT 2.260 1.445 2.565 1.615 ;
        RECT 2.260 1.245 2.430 1.445 ;
        RECT 1.875 1.075 2.430 1.245 ;
        RECT 2.215 0.895 2.430 1.075 ;
        RECT 0.085 0.085 0.365 0.895 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.895 ;
        RECT 2.215 0.725 2.565 0.895 ;
        RECT 2.395 0.445 2.565 0.725 ;
        RECT 2.775 0.085 3.030 0.845 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_2

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_isobufsrc_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.075 4.975 1.320 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.360 1.075 1.800 1.275 ;
    END
  END SLEEP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.875 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER li1 ;
        RECT 2.295 1.745 2.465 2.125 ;
        RECT 3.135 1.745 3.305 2.125 ;
        RECT 2.295 1.445 3.305 1.745 ;
        RECT 2.295 0.905 2.625 1.445 ;
        RECT 0.535 0.725 3.385 0.905 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 3.055 0.255 3.385 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.085 1.665 0.365 2.465 ;
        RECT 0.535 1.835 0.865 2.635 ;
        RECT 1.035 1.665 1.205 2.465 ;
        RECT 1.375 1.835 1.625 2.635 ;
        RECT 1.795 2.295 3.855 2.465 ;
        RECT 1.795 1.665 2.125 2.295 ;
        RECT 2.635 1.935 2.965 2.295 ;
        RECT 0.085 1.455 2.125 1.665 ;
        RECT 3.475 1.575 3.855 2.295 ;
        RECT 4.025 1.575 4.355 2.465 ;
        RECT 4.025 1.275 4.275 1.575 ;
        RECT 4.525 1.495 4.930 2.635 ;
        RECT 2.795 1.075 4.275 1.275 ;
        RECT 0.085 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.555 ;
        RECT 2.715 0.085 2.885 0.555 ;
        RECT 3.555 0.085 3.845 0.905 ;
        RECT 4.025 0.815 4.275 1.075 ;
        RECT 4.025 0.255 4.355 0.815 ;
        RECT 4.525 0.085 4.815 0.905 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_4

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_isobufsrc_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.065 0.575 1.285 ;
        RECT 0.085 0.255 0.265 1.065 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 5.270 1.075 8.010 1.275 ;
    END
  END SLEEP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484000 ;
    PORT
      LAYER li1 ;
        RECT 5.405 1.615 5.655 2.125 ;
        RECT 6.245 1.615 6.495 2.125 ;
        RECT 7.085 1.615 7.335 2.125 ;
        RECT 7.925 1.615 8.175 2.125 ;
        RECT 5.405 1.445 8.655 1.615 ;
        RECT 8.180 0.905 8.655 1.445 ;
        RECT 2.005 0.725 8.655 0.905 ;
        RECT 2.005 0.255 2.335 0.725 ;
        RECT 2.845 0.255 3.175 0.725 ;
        RECT 3.685 0.255 4.015 0.725 ;
        RECT 4.525 0.255 4.855 0.725 ;
        RECT 5.365 0.255 5.695 0.725 ;
        RECT 6.205 0.255 6.535 0.725 ;
        RECT 7.045 0.255 7.375 0.725 ;
        RECT 7.885 0.255 8.215 0.725 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 0.315 0.105 8.725 1.015 ;
      LAYER li1 ;
        RECT 0.000 2.635 8.740 2.805 ;
        RECT 0.195 1.455 0.415 2.635 ;
        RECT 0.585 1.455 0.915 2.465 ;
        RECT 1.085 1.455 1.330 2.635 ;
        RECT 1.555 1.665 1.875 2.465 ;
        RECT 2.045 1.835 2.295 2.635 ;
        RECT 2.465 1.665 2.715 2.465 ;
        RECT 2.885 1.835 3.135 2.635 ;
        RECT 3.305 1.665 3.555 2.465 ;
        RECT 3.725 1.835 3.975 2.635 ;
        RECT 4.145 1.665 4.395 2.465 ;
        RECT 4.565 1.835 4.815 2.635 ;
        RECT 4.985 2.295 8.595 2.465 ;
        RECT 4.985 1.665 5.235 2.295 ;
        RECT 5.825 1.785 6.075 2.295 ;
        RECT 6.665 1.785 6.915 2.295 ;
        RECT 7.505 1.785 7.755 2.295 ;
        RECT 8.345 1.785 8.595 2.295 ;
        RECT 1.555 1.455 5.235 1.665 ;
        RECT 0.745 1.285 0.915 1.455 ;
        RECT 0.745 1.075 5.000 1.285 ;
        RECT 0.745 1.065 1.155 1.075 ;
        RECT 0.435 0.085 0.655 0.895 ;
        RECT 0.825 0.255 1.155 1.065 ;
        RECT 1.325 0.085 1.835 0.905 ;
        RECT 2.505 0.085 2.675 0.555 ;
        RECT 3.345 0.085 3.515 0.555 ;
        RECT 4.185 0.085 4.355 0.555 ;
        RECT 5.025 0.085 5.195 0.555 ;
        RECT 5.865 0.085 6.035 0.555 ;
        RECT 6.705 0.085 6.875 0.555 ;
        RECT 7.545 0.085 7.715 0.555 ;
        RECT 8.385 0.085 8.655 0.555 ;
        RECT 0.000 -0.085 8.740 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_8

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_isobufsrc_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrc_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.560 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.665 1.325 ;
        RECT 0.085 0.255 0.315 0.995 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.960000 ;
    PORT
      LAYER li1 ;
        RECT 9.450 1.075 15.650 1.285 ;
    END
  END SLEEP
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 16.560 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 16.750 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 16.560 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.968000 ;
    PORT
      LAYER li1 ;
        RECT 9.685 1.625 9.935 2.125 ;
        RECT 10.525 1.625 10.775 2.125 ;
        RECT 11.365 1.625 11.615 2.125 ;
        RECT 12.205 1.625 12.455 2.125 ;
        RECT 13.045 1.625 13.295 2.125 ;
        RECT 13.885 1.625 14.135 2.125 ;
        RECT 14.725 1.625 14.975 2.125 ;
        RECT 15.565 1.625 15.815 2.125 ;
        RECT 9.685 1.455 16.475 1.625 ;
        RECT 15.820 0.905 16.475 1.455 ;
        RECT 2.925 0.725 16.475 0.905 ;
        RECT 2.925 0.255 3.255 0.725 ;
        RECT 3.765 0.255 4.095 0.725 ;
        RECT 4.605 0.255 4.935 0.725 ;
        RECT 5.445 0.255 5.775 0.725 ;
        RECT 6.285 0.255 6.615 0.725 ;
        RECT 7.125 0.255 7.455 0.725 ;
        RECT 7.965 0.255 8.295 0.725 ;
        RECT 8.805 0.255 9.135 0.725 ;
        RECT 9.645 0.255 9.975 0.725 ;
        RECT 10.485 0.255 10.815 0.725 ;
        RECT 11.325 0.255 11.655 0.725 ;
        RECT 12.165 0.255 12.495 0.725 ;
        RECT 13.005 0.255 13.335 0.725 ;
        RECT 13.845 0.255 14.175 0.725 ;
        RECT 14.685 0.255 15.015 0.725 ;
        RECT 15.525 0.255 15.855 0.725 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 0.395 0.105 16.365 1.015 ;
      LAYER li1 ;
        RECT 0.000 2.635 16.560 2.805 ;
        RECT 0.300 1.495 0.515 2.635 ;
        RECT 0.685 1.495 1.015 2.465 ;
        RECT 0.835 1.285 1.015 1.495 ;
        RECT 1.185 1.455 1.355 2.635 ;
        RECT 1.525 1.285 1.855 2.465 ;
        RECT 2.025 1.455 2.270 2.635 ;
        RECT 2.475 1.665 2.795 2.465 ;
        RECT 2.965 1.835 3.215 2.635 ;
        RECT 3.385 1.665 3.635 2.465 ;
        RECT 3.805 1.835 4.055 2.635 ;
        RECT 4.225 1.665 4.475 2.465 ;
        RECT 4.645 1.835 4.895 2.635 ;
        RECT 5.065 1.665 5.315 2.465 ;
        RECT 5.485 1.835 5.735 2.635 ;
        RECT 5.905 1.665 6.155 2.465 ;
        RECT 6.325 1.835 6.575 2.635 ;
        RECT 6.745 1.665 6.995 2.465 ;
        RECT 7.165 1.835 7.415 2.635 ;
        RECT 7.585 1.665 7.835 2.465 ;
        RECT 8.005 1.835 8.255 2.635 ;
        RECT 8.425 1.665 8.675 2.465 ;
        RECT 8.845 1.835 9.095 2.635 ;
        RECT 9.265 2.295 16.235 2.465 ;
        RECT 9.265 1.665 9.515 2.295 ;
        RECT 10.105 1.795 10.355 2.295 ;
        RECT 10.945 1.795 11.195 2.295 ;
        RECT 11.785 1.795 12.035 2.295 ;
        RECT 12.625 1.795 12.875 2.295 ;
        RECT 13.465 1.795 13.715 2.295 ;
        RECT 14.305 1.795 14.555 2.295 ;
        RECT 15.145 1.795 15.395 2.295 ;
        RECT 15.985 1.795 16.235 2.295 ;
        RECT 2.475 1.455 9.515 1.665 ;
        RECT 0.835 1.075 9.280 1.285 ;
        RECT 0.835 1.065 2.035 1.075 ;
        RECT 0.485 0.085 0.815 0.825 ;
        RECT 0.985 0.255 1.195 1.065 ;
        RECT 1.365 0.085 1.615 0.895 ;
        RECT 1.785 0.255 2.035 1.065 ;
        RECT 2.205 0.085 2.755 0.905 ;
        RECT 3.425 0.085 3.595 0.555 ;
        RECT 4.265 0.085 4.435 0.555 ;
        RECT 5.105 0.085 5.275 0.555 ;
        RECT 5.945 0.085 6.115 0.555 ;
        RECT 6.785 0.085 6.955 0.555 ;
        RECT 7.625 0.085 7.795 0.555 ;
        RECT 8.465 0.085 8.635 0.555 ;
        RECT 9.305 0.085 9.475 0.555 ;
        RECT 10.145 0.085 10.315 0.555 ;
        RECT 10.985 0.085 11.155 0.555 ;
        RECT 11.825 0.085 11.995 0.555 ;
        RECT 12.665 0.085 12.835 0.555 ;
        RECT 13.505 0.085 13.675 0.555 ;
        RECT 14.345 0.085 14.515 0.555 ;
        RECT 15.185 0.085 15.355 0.555 ;
        RECT 16.025 0.085 16.295 0.555 ;
        RECT 0.000 -0.085 16.560 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 15.325 2.635 15.495 2.805 ;
        RECT 15.785 2.635 15.955 2.805 ;
        RECT 16.245 2.635 16.415 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
        RECT 15.325 -0.085 15.495 0.085 ;
        RECT 15.785 -0.085 15.955 0.085 ;
        RECT 16.245 -0.085 16.415 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrc_16

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_isobufsrckapwr_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.260 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.615 1.320 ;
    END
  END A
  PIN SLEEP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.260 1.075 4.700 1.275 ;
    END
  END SLEEP
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.070 2.140 14.190 2.340 ;
        RECT 5.175 2.080 5.465 2.140 ;
        RECT 6.035 2.080 6.325 2.140 ;
        RECT 6.890 2.080 7.180 2.140 ;
        RECT 7.740 2.080 8.030 2.140 ;
        RECT 8.620 2.080 8.910 2.140 ;
        RECT 9.480 2.080 9.770 2.140 ;
        RECT 10.335 2.080 10.625 2.140 ;
        RECT 11.195 2.080 11.485 2.140 ;
        RECT 12.050 2.080 12.340 2.140 ;
        RECT 12.900 2.080 13.190 2.140 ;
        RECT 13.780 2.080 14.070 2.140 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 14.260 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.185 0.785 5.055 1.015 ;
        RECT 0.185 0.105 14.170 0.785 ;
        RECT 0.185 0.085 0.320 0.105 ;
        RECT 0.150 -0.085 0.320 0.085 ;
        RECT 5.205 -0.085 5.375 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 14.450 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 14.260 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER li1 ;
        RECT 7.375 1.735 7.600 2.460 ;
        RECT 8.200 1.735 8.460 2.460 ;
        RECT 9.060 1.735 9.320 2.460 ;
        RECT 9.920 1.735 10.180 2.460 ;
        RECT 10.765 1.735 11.025 2.460 ;
        RECT 11.625 1.735 11.885 2.460 ;
        RECT 12.485 1.735 12.745 2.460 ;
        RECT 7.375 1.720 12.745 1.735 ;
        RECT 13.355 1.720 13.645 2.460 ;
        RECT 7.375 1.495 14.085 1.720 ;
        RECT 12.920 0.905 14.085 1.495 ;
        RECT 7.340 0.735 14.085 0.905 ;
        RECT 7.340 0.280 7.600 0.735 ;
        RECT 8.200 0.280 8.460 0.735 ;
        RECT 9.060 0.280 9.320 0.735 ;
        RECT 9.905 0.280 10.180 0.735 ;
        RECT 10.765 0.280 11.025 0.735 ;
        RECT 11.625 0.280 11.885 0.735 ;
        RECT 12.485 0.280 12.745 0.735 ;
        RECT 13.355 0.280 13.615 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 14.260 2.805 ;
        RECT 0.130 1.495 0.535 2.635 ;
        RECT 0.705 1.575 1.035 2.465 ;
        RECT 1.205 2.295 3.265 2.465 ;
        RECT 1.205 1.575 1.585 2.295 ;
        RECT 1.755 1.745 1.925 2.125 ;
        RECT 2.095 1.935 2.425 2.295 ;
        RECT 2.595 1.745 2.765 2.125 ;
        RECT 0.785 1.275 1.035 1.575 ;
        RECT 1.755 1.445 2.765 1.745 ;
        RECT 2.935 1.665 3.265 2.295 ;
        RECT 3.435 1.835 3.685 2.635 ;
        RECT 3.855 1.665 4.025 2.465 ;
        RECT 4.195 1.835 4.525 2.635 ;
        RECT 4.695 1.665 4.975 2.465 ;
        RECT 2.935 1.455 4.975 1.665 ;
        RECT 5.155 1.495 5.485 2.465 ;
        RECT 0.785 1.075 2.265 1.275 ;
        RECT 0.245 0.085 0.535 0.905 ;
        RECT 0.785 0.815 1.035 1.075 ;
        RECT 2.435 0.965 2.765 1.445 ;
        RECT 5.655 1.325 5.845 2.465 ;
        RECT 6.015 1.495 6.345 2.465 ;
        RECT 6.515 1.325 6.705 2.460 ;
        RECT 6.875 1.495 7.205 2.465 ;
        RECT 7.770 1.905 8.030 2.465 ;
        RECT 8.630 1.905 8.890 2.465 ;
        RECT 9.490 1.905 9.750 2.465 ;
        RECT 10.350 1.905 10.595 2.465 ;
        RECT 11.210 1.905 11.455 2.465 ;
        RECT 12.070 1.905 12.315 2.465 ;
        RECT 12.930 1.905 13.185 2.465 ;
        RECT 13.815 1.890 14.085 2.465 ;
        RECT 2.435 0.905 3.095 0.965 ;
        RECT 0.705 0.255 1.035 0.815 ;
        RECT 1.215 0.085 1.505 0.905 ;
        RECT 1.675 0.725 4.525 0.905 ;
        RECT 1.675 0.255 2.005 0.725 ;
        RECT 2.175 0.085 2.345 0.555 ;
        RECT 2.515 0.255 2.845 0.725 ;
        RECT 3.015 0.085 3.185 0.555 ;
        RECT 3.355 0.255 3.685 0.725 ;
        RECT 3.855 0.085 4.025 0.555 ;
        RECT 4.195 0.255 4.525 0.725 ;
        RECT 4.695 0.565 4.975 0.905 ;
        RECT 5.145 0.735 5.460 1.325 ;
        RECT 5.655 1.075 12.750 1.325 ;
        RECT 4.695 0.085 5.450 0.565 ;
        RECT 5.655 0.265 5.880 1.075 ;
        RECT 6.050 0.085 6.310 0.610 ;
        RECT 6.490 0.265 6.740 1.075 ;
        RECT 6.910 0.085 7.170 0.645 ;
        RECT 7.770 0.085 8.030 0.565 ;
        RECT 8.630 0.085 8.890 0.565 ;
        RECT 9.490 0.085 9.735 0.565 ;
        RECT 10.350 0.085 10.595 0.565 ;
        RECT 11.205 0.085 11.455 0.565 ;
        RECT 12.065 0.085 12.315 0.565 ;
        RECT 12.925 0.085 13.185 0.565 ;
        RECT 13.785 0.085 14.085 0.565 ;
        RECT 0.000 -0.085 14.260 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 5.235 2.125 5.405 2.295 ;
        RECT 6.095 2.125 6.265 2.295 ;
        RECT 6.950 2.125 7.120 2.295 ;
        RECT 7.800 2.125 7.970 2.295 ;
        RECT 8.680 2.125 8.850 2.295 ;
        RECT 9.540 2.125 9.710 2.295 ;
        RECT 10.395 2.125 10.565 2.295 ;
        RECT 11.255 2.125 11.425 2.295 ;
        RECT 12.110 2.125 12.280 2.295 ;
        RECT 12.960 2.125 13.130 2.295 ;
        RECT 13.840 2.125 14.010 2.295 ;
        RECT 2.525 0.765 2.695 0.935 ;
        RECT 2.885 0.765 3.055 0.935 ;
        RECT 5.210 0.765 5.380 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
      LAYER met1 ;
        RECT 2.465 0.920 3.115 0.965 ;
        RECT 5.150 0.920 5.440 0.965 ;
        RECT 2.465 0.780 5.440 0.920 ;
        RECT 2.465 0.735 3.115 0.780 ;
        RECT 5.150 0.735 5.440 0.780 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrckapwr_16

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 5.440 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.603000 ;
    PORT
      LAYER li1 ;
        RECT 2.970 1.070 3.290 1.540 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 2.555 5.250 5.555 5.335 ;
        RECT 0.015 4.465 0.445 5.250 ;
        RECT 2.555 4.465 6.225 5.250 ;
        RECT 2.555 4.425 5.555 4.465 ;
      LAYER met1 ;
        RECT 0.000 5.200 6.440 5.680 ;
    END
    PORT
      LAYER pwell ;
        RECT 3.005 0.975 5.705 1.070 ;
        RECT 0.015 0.190 0.445 0.975 ;
        RECT 3.005 0.960 6.225 0.975 ;
        RECT 1.990 0.280 6.225 0.960 ;
        RECT 3.005 0.190 6.225 0.280 ;
        RECT 3.005 0.160 5.705 0.190 ;
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 4.135 ;
        RECT 4.250 1.305 6.630 4.135 ;
      LAYER met1 ;
        RECT 0.080 3.640 0.370 3.685 ;
        RECT 5.870 3.640 6.160 3.685 ;
        RECT 0.070 3.500 6.170 3.640 ;
        RECT 0.080 3.455 0.370 3.500 ;
        RECT 5.870 3.455 6.160 3.500 ;
    END
  END VPB
  PIN VPWRIN
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 1.920 1.305 2.980 4.135 ;
      LAYER met1 ;
        RECT 1.360 2.280 2.370 2.315 ;
        RECT 0.070 2.140 6.170 2.280 ;
        RECT 1.360 2.085 2.370 2.140 ;
    END
  END VPWRIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.402500 ;
    PORT
      LAYER li1 ;
        RECT 5.360 0.980 5.635 2.370 ;
        RECT 5.335 0.290 5.635 0.980 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 5.355 6.440 5.525 ;
        RECT 0.085 4.630 0.375 5.355 ;
        RECT 2.645 4.515 2.905 5.355 ;
        RECT 3.075 4.325 3.405 5.185 ;
        RECT 3.575 4.515 3.765 5.355 ;
        RECT 3.935 4.325 4.265 5.185 ;
        RECT 4.445 4.515 4.955 5.355 ;
        RECT 5.135 4.820 5.485 5.160 ;
        RECT 5.135 4.460 5.695 4.820 ;
        RECT 5.865 4.630 6.155 5.355 ;
        RECT 5.135 4.405 5.765 4.460 ;
        RECT 3.075 4.265 4.265 4.325 ;
        RECT 5.360 4.355 5.765 4.405 ;
        RECT 3.145 4.155 4.195 4.265 ;
        RECT 0.085 2.985 0.375 3.970 ;
        RECT 0.000 2.635 1.890 2.805 ;
        RECT 2.060 2.660 2.810 3.750 ;
        RECT 2.060 2.335 2.390 2.660 ;
        RECT 3.060 2.370 3.390 3.965 ;
        RECT 4.020 3.810 4.190 4.155 ;
        RECT 5.360 4.125 6.085 4.355 ;
        RECT 4.410 3.640 4.720 3.740 ;
        RECT 3.680 3.470 4.720 3.640 ;
        RECT 3.680 2.575 3.850 3.470 ;
        RECT 4.020 2.915 4.190 3.300 ;
        RECT 4.390 3.085 4.720 3.470 ;
        RECT 4.020 2.745 4.640 2.915 ;
        RECT 3.680 2.405 4.190 2.575 ;
        RECT 1.380 2.065 2.390 2.335 ;
        RECT 2.060 1.635 2.390 2.065 ;
        RECT 2.560 2.130 3.390 2.370 ;
        RECT 0.085 0.085 0.375 0.810 ;
        RECT 2.020 0.085 2.350 0.895 ;
        RECT 2.560 0.375 2.800 2.130 ;
        RECT 4.020 0.980 4.190 2.405 ;
        RECT 4.470 1.625 4.640 2.745 ;
        RECT 4.890 2.805 5.120 3.740 ;
        RECT 5.360 3.070 5.550 4.125 ;
        RECT 5.865 2.985 6.155 3.955 ;
        RECT 4.890 2.635 6.440 2.805 ;
        RECT 4.890 1.625 5.120 2.635 ;
        RECT 3.115 0.085 3.445 0.900 ;
        RECT 3.615 0.730 4.665 0.980 ;
        RECT 3.615 0.290 3.805 0.730 ;
        RECT 3.975 0.085 4.305 0.560 ;
        RECT 4.475 0.290 4.665 0.730 ;
        RECT 4.835 0.085 5.165 0.900 ;
        RECT 5.865 0.085 6.155 0.810 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 5.355 0.315 5.525 ;
        RECT 0.605 5.355 0.775 5.525 ;
        RECT 1.065 5.355 1.235 5.525 ;
        RECT 1.525 5.355 1.695 5.525 ;
        RECT 1.985 5.355 2.155 5.525 ;
        RECT 2.445 5.355 2.615 5.525 ;
        RECT 2.905 5.355 3.075 5.525 ;
        RECT 3.365 5.355 3.535 5.525 ;
        RECT 3.825 5.355 3.995 5.525 ;
        RECT 4.285 5.355 4.455 5.525 ;
        RECT 4.745 5.355 4.915 5.525 ;
        RECT 5.205 5.355 5.375 5.525 ;
        RECT 5.665 5.355 5.835 5.525 ;
        RECT 6.125 5.355 6.295 5.525 ;
        RECT 0.140 3.485 0.310 3.655 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.420 2.115 1.590 2.285 ;
        RECT 1.780 2.115 1.950 2.285 ;
        RECT 2.140 2.115 2.310 2.285 ;
        RECT 5.930 3.485 6.100 3.655 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_1

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 5.440 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.603000 ;
    PORT
      LAYER li1 ;
        RECT 2.970 1.070 3.290 1.540 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 2.555 5.250 5.555 5.335 ;
        RECT 0.015 4.465 0.445 5.250 ;
        RECT 2.555 4.465 6.425 5.250 ;
        RECT 2.555 4.425 5.555 4.465 ;
      LAYER met1 ;
        RECT 0.000 5.200 6.440 5.680 ;
    END
    PORT
      LAYER pwell ;
        RECT 0.015 0.190 0.445 0.975 ;
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 4.135 ;
        RECT 4.250 1.305 6.630 4.135 ;
      LAYER met1 ;
        RECT 0.080 3.640 0.370 3.685 ;
        RECT 6.010 3.640 6.300 3.685 ;
        RECT 0.070 3.500 6.300 3.640 ;
        RECT 0.080 3.455 0.370 3.500 ;
        RECT 6.010 3.455 6.300 3.500 ;
    END
  END VPB
  PIN VPWRIN
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 1.920 1.305 2.980 4.135 ;
      LAYER met1 ;
        RECT 1.360 2.280 2.370 2.315 ;
        RECT 0.070 2.140 6.370 2.280 ;
        RECT 1.360 2.085 2.370 2.140 ;
    END
  END VPWRIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.610500 ;
    PORT
      LAYER li1 ;
        RECT 5.360 0.980 5.635 2.370 ;
        RECT 5.335 0.255 5.635 0.980 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 3.005 0.960 6.265 1.015 ;
        RECT 1.990 0.280 6.265 0.960 ;
        RECT 3.005 0.105 6.265 0.280 ;
      LAYER li1 ;
        RECT 0.000 5.355 6.440 5.525 ;
        RECT 0.085 4.630 0.375 5.355 ;
        RECT 2.645 4.515 2.905 5.355 ;
        RECT 3.075 4.325 3.405 5.185 ;
        RECT 3.575 4.515 3.765 5.355 ;
        RECT 3.935 4.325 4.265 5.185 ;
        RECT 4.445 4.515 4.955 5.355 ;
        RECT 5.135 4.820 5.485 5.160 ;
        RECT 5.135 4.460 5.695 4.820 ;
        RECT 6.065 4.630 6.355 5.355 ;
        RECT 5.135 4.405 5.765 4.460 ;
        RECT 3.075 4.265 4.265 4.325 ;
        RECT 5.360 4.355 5.765 4.405 ;
        RECT 3.145 4.155 4.195 4.265 ;
        RECT 0.085 2.985 0.375 3.970 ;
        RECT 0.000 2.635 1.890 2.805 ;
        RECT 2.060 2.660 2.810 3.750 ;
        RECT 2.060 2.335 2.390 2.660 ;
        RECT 3.060 2.370 3.390 3.965 ;
        RECT 4.020 3.810 4.190 4.155 ;
        RECT 5.360 4.125 6.085 4.355 ;
        RECT 4.410 3.640 4.720 3.740 ;
        RECT 3.680 3.470 4.720 3.640 ;
        RECT 3.680 2.575 3.850 3.470 ;
        RECT 4.020 2.915 4.190 3.300 ;
        RECT 4.390 3.085 4.720 3.470 ;
        RECT 4.020 2.745 4.640 2.915 ;
        RECT 3.680 2.405 4.190 2.575 ;
        RECT 1.380 2.065 2.390 2.335 ;
        RECT 2.060 1.635 2.390 2.065 ;
        RECT 2.560 2.130 3.390 2.370 ;
        RECT 0.085 0.085 0.375 0.810 ;
        RECT 2.020 0.085 2.350 0.895 ;
        RECT 2.560 0.375 2.800 2.130 ;
        RECT 4.020 0.980 4.190 2.405 ;
        RECT 4.470 1.625 4.640 2.745 ;
        RECT 4.890 2.805 5.120 3.740 ;
        RECT 5.360 3.070 5.550 4.125 ;
        RECT 6.065 2.985 6.355 3.955 ;
        RECT 4.890 2.635 6.440 2.805 ;
        RECT 4.890 1.625 5.120 2.635 ;
        RECT 5.905 1.610 6.075 2.635 ;
        RECT 3.115 0.085 3.445 0.900 ;
        RECT 3.615 0.730 4.665 0.980 ;
        RECT 3.615 0.255 3.805 0.730 ;
        RECT 3.975 0.085 4.305 0.560 ;
        RECT 4.475 0.255 4.665 0.730 ;
        RECT 4.835 0.085 5.165 0.900 ;
        RECT 5.825 0.085 6.155 0.900 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 5.355 0.315 5.525 ;
        RECT 0.605 5.355 0.775 5.525 ;
        RECT 1.065 5.355 1.235 5.525 ;
        RECT 1.525 5.355 1.695 5.525 ;
        RECT 1.985 5.355 2.155 5.525 ;
        RECT 2.445 5.355 2.615 5.525 ;
        RECT 2.905 5.355 3.075 5.525 ;
        RECT 3.365 5.355 3.535 5.525 ;
        RECT 3.825 5.355 3.995 5.525 ;
        RECT 4.285 5.355 4.455 5.525 ;
        RECT 4.745 5.355 4.915 5.525 ;
        RECT 5.205 5.355 5.375 5.525 ;
        RECT 5.665 5.355 5.835 5.525 ;
        RECT 6.125 5.355 6.295 5.525 ;
        RECT 0.140 3.485 0.310 3.655 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.420 2.115 1.590 2.285 ;
        RECT 1.780 2.115 1.950 2.285 ;
        RECT 2.140 2.115 2.310 2.285 ;
        RECT 6.070 3.485 6.240 3.655 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_2

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 5.440 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.603000 ;
    PORT
      LAYER li1 ;
        RECT 2.970 1.070 3.290 1.540 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 0.015 4.465 0.445 5.250 ;
        RECT 6.915 4.465 7.345 5.250 ;
      LAYER met1 ;
        RECT 0.000 5.200 7.360 5.680 ;
    END
    PORT
      LAYER pwell ;
        RECT 0.015 0.190 0.445 0.975 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 4.135 ;
        RECT 4.250 1.305 7.405 4.135 ;
      LAYER met1 ;
        RECT 0.080 3.640 0.370 3.685 ;
        RECT 6.930 3.640 7.220 3.685 ;
        RECT 0.070 3.500 7.290 3.640 ;
        RECT 0.080 3.455 0.370 3.500 ;
        RECT 6.930 3.455 7.220 3.500 ;
    END
  END VPB
  PIN VPWRIN
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 1.920 1.305 2.980 4.135 ;
      LAYER met1 ;
        RECT 1.360 2.280 2.370 2.315 ;
        RECT 0.070 2.140 7.290 2.280 ;
        RECT 1.360 2.085 2.370 2.140 ;
    END
  END VPWRIN
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.072500 ;
    PORT
      LAYER li1 ;
        RECT 5.360 1.410 5.635 2.370 ;
        RECT 6.280 1.410 6.555 2.370 ;
        RECT 5.360 1.085 6.555 1.410 ;
        RECT 5.360 0.980 5.635 1.085 ;
        RECT 5.335 0.255 5.635 0.980 ;
        RECT 6.335 0.255 6.555 1.085 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 2.555 4.425 5.555 5.335 ;
        RECT 3.005 0.960 7.125 1.015 ;
        RECT 1.990 0.280 7.125 0.960 ;
        RECT 3.005 0.105 7.125 0.280 ;
      LAYER li1 ;
        RECT 0.000 5.355 7.360 5.525 ;
        RECT 0.085 4.630 0.375 5.355 ;
        RECT 2.645 4.515 2.905 5.355 ;
        RECT 3.075 4.325 3.405 5.185 ;
        RECT 3.575 4.515 3.765 5.355 ;
        RECT 3.935 4.325 4.265 5.185 ;
        RECT 4.445 4.515 4.955 5.355 ;
        RECT 5.135 4.820 5.485 5.160 ;
        RECT 5.135 4.460 5.695 4.820 ;
        RECT 6.985 4.630 7.275 5.355 ;
        RECT 5.135 4.405 5.765 4.460 ;
        RECT 3.075 4.265 4.265 4.325 ;
        RECT 5.360 4.355 5.765 4.405 ;
        RECT 3.145 4.155 4.195 4.265 ;
        RECT 0.085 2.985 0.375 3.970 ;
        RECT 0.000 2.635 1.890 2.805 ;
        RECT 2.060 2.660 2.810 3.750 ;
        RECT 2.060 2.335 2.390 2.660 ;
        RECT 3.060 2.370 3.390 3.965 ;
        RECT 4.020 3.810 4.190 4.155 ;
        RECT 5.360 4.125 6.085 4.355 ;
        RECT 4.410 3.640 4.720 3.740 ;
        RECT 3.680 3.470 4.720 3.640 ;
        RECT 3.680 2.575 3.850 3.470 ;
        RECT 4.020 2.915 4.190 3.300 ;
        RECT 4.390 3.085 4.720 3.470 ;
        RECT 4.020 2.745 4.640 2.915 ;
        RECT 3.680 2.405 4.190 2.575 ;
        RECT 1.380 2.065 2.390 2.335 ;
        RECT 2.060 1.635 2.390 2.065 ;
        RECT 2.560 2.130 3.390 2.370 ;
        RECT 0.085 0.085 0.375 0.810 ;
        RECT 2.020 0.085 2.350 0.895 ;
        RECT 2.560 0.375 2.800 2.130 ;
        RECT 4.020 0.980 4.190 2.405 ;
        RECT 4.470 1.625 4.640 2.745 ;
        RECT 4.890 2.805 5.120 3.740 ;
        RECT 5.360 3.070 5.550 4.125 ;
        RECT 6.985 2.985 7.275 3.955 ;
        RECT 4.890 2.635 7.360 2.805 ;
        RECT 4.890 1.625 5.120 2.635 ;
        RECT 5.905 1.610 6.075 2.635 ;
        RECT 6.755 1.610 6.935 2.635 ;
        RECT 3.115 0.085 3.445 0.900 ;
        RECT 3.615 0.730 4.665 0.980 ;
        RECT 3.615 0.255 3.805 0.730 ;
        RECT 3.975 0.085 4.305 0.560 ;
        RECT 4.475 0.255 4.665 0.730 ;
        RECT 4.835 0.085 5.165 0.900 ;
        RECT 5.825 0.085 6.155 0.845 ;
        RECT 6.755 0.085 7.005 0.925 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 5.355 0.315 5.525 ;
        RECT 0.605 5.355 0.775 5.525 ;
        RECT 1.065 5.355 1.235 5.525 ;
        RECT 1.525 5.355 1.695 5.525 ;
        RECT 1.985 5.355 2.155 5.525 ;
        RECT 2.445 5.355 2.615 5.525 ;
        RECT 2.905 5.355 3.075 5.525 ;
        RECT 3.365 5.355 3.535 5.525 ;
        RECT 3.825 5.355 3.995 5.525 ;
        RECT 4.285 5.355 4.455 5.525 ;
        RECT 4.745 5.355 4.915 5.525 ;
        RECT 5.205 5.355 5.375 5.525 ;
        RECT 5.665 5.355 5.835 5.525 ;
        RECT 6.125 5.355 6.295 5.525 ;
        RECT 6.585 5.355 6.755 5.525 ;
        RECT 7.045 5.355 7.215 5.525 ;
        RECT 0.140 3.485 0.310 3.655 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.420 2.115 1.590 2.285 ;
        RECT 1.780 2.115 1.950 2.285 ;
        RECT 2.140 2.115 2.310 2.285 ;
        RECT 6.990 3.485 7.160 3.655 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_hl_isowell_tap_4

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 5.440 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.603000 ;
    PORT
      LAYER li1 ;
        RECT 2.970 1.070 3.290 1.540 ;
    END
  END A
  PIN LOWLVPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 1.920 1.305 2.980 4.135 ;
      LAYER met1 ;
        RECT 1.360 2.280 2.370 2.315 ;
        RECT 0.070 2.140 7.290 2.280 ;
        RECT 1.360 2.085 2.370 2.140 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 5.200 7.360 5.680 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.075 5.245 0.200 5.395 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 4.250 1.305 7.405 4.135 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.072500 ;
    PORT
      LAYER li1 ;
        RECT 5.360 1.410 5.635 2.370 ;
        RECT 6.280 1.410 6.555 2.370 ;
        RECT 5.360 1.085 6.555 1.410 ;
        RECT 5.360 0.980 5.635 1.085 ;
        RECT 5.335 0.255 5.635 0.980 ;
        RECT 6.335 0.255 6.555 1.085 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 2.555 4.425 5.555 5.335 ;
      LAYER nwell ;
        RECT -0.190 1.305 0.650 4.135 ;
      LAYER pwell ;
        RECT 3.005 0.960 7.125 1.015 ;
        RECT 1.990 0.280 7.125 0.960 ;
        RECT 3.005 0.105 7.125 0.280 ;
      LAYER li1 ;
        RECT 0.000 5.355 7.360 5.525 ;
        RECT 2.645 4.515 2.905 5.355 ;
        RECT 3.075 4.325 3.405 5.185 ;
        RECT 3.575 4.515 3.765 5.355 ;
        RECT 3.935 4.325 4.265 5.185 ;
        RECT 4.445 4.515 4.955 5.355 ;
        RECT 5.135 4.820 5.485 5.160 ;
        RECT 5.135 4.460 5.695 4.820 ;
        RECT 5.135 4.405 5.765 4.460 ;
        RECT 3.075 4.265 4.265 4.325 ;
        RECT 5.360 4.355 5.765 4.405 ;
        RECT 3.145 4.155 4.195 4.265 ;
        RECT 0.000 2.635 1.890 2.805 ;
        RECT 2.060 2.660 2.810 3.750 ;
        RECT 2.060 2.335 2.390 2.660 ;
        RECT 3.060 2.370 3.390 3.965 ;
        RECT 4.020 3.810 4.190 4.155 ;
        RECT 5.360 4.125 6.085 4.355 ;
        RECT 4.410 3.640 4.720 3.740 ;
        RECT 3.680 3.470 4.720 3.640 ;
        RECT 3.680 2.575 3.850 3.470 ;
        RECT 4.020 2.915 4.190 3.300 ;
        RECT 4.390 3.085 4.720 3.470 ;
        RECT 4.020 2.745 4.640 2.915 ;
        RECT 3.680 2.405 4.190 2.575 ;
        RECT 1.380 2.065 2.390 2.335 ;
        RECT 2.060 1.635 2.390 2.065 ;
        RECT 2.560 2.130 3.390 2.370 ;
        RECT 2.020 0.085 2.350 0.895 ;
        RECT 2.560 0.375 2.800 2.130 ;
        RECT 4.020 0.980 4.190 2.405 ;
        RECT 4.470 1.625 4.640 2.745 ;
        RECT 4.890 2.805 5.120 3.740 ;
        RECT 5.360 3.070 5.550 4.125 ;
        RECT 4.890 2.635 7.360 2.805 ;
        RECT 4.890 1.625 5.120 2.635 ;
        RECT 5.905 1.610 6.075 2.635 ;
        RECT 6.755 1.610 6.935 2.635 ;
        RECT 3.115 0.085 3.445 0.900 ;
        RECT 3.615 0.730 4.665 0.980 ;
        RECT 3.615 0.255 3.805 0.730 ;
        RECT 3.975 0.085 4.305 0.560 ;
        RECT 4.475 0.255 4.665 0.730 ;
        RECT 4.835 0.085 5.165 0.900 ;
        RECT 5.825 0.085 6.155 0.845 ;
        RECT 6.755 0.085 7.005 0.925 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 5.355 0.315 5.525 ;
        RECT 0.605 5.355 0.775 5.525 ;
        RECT 1.065 5.355 1.235 5.525 ;
        RECT 1.525 5.355 1.695 5.525 ;
        RECT 1.985 5.355 2.155 5.525 ;
        RECT 2.445 5.355 2.615 5.525 ;
        RECT 2.905 5.355 3.075 5.525 ;
        RECT 3.365 5.355 3.535 5.525 ;
        RECT 3.825 5.355 3.995 5.525 ;
        RECT 4.285 5.355 4.455 5.525 ;
        RECT 4.745 5.355 4.915 5.525 ;
        RECT 5.205 5.355 5.375 5.525 ;
        RECT 5.665 5.355 5.835 5.525 ;
        RECT 6.125 5.355 6.295 5.525 ;
        RECT 6.585 5.355 6.755 5.525 ;
        RECT 7.045 5.355 7.215 5.525 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.420 2.115 1.590 2.285 ;
        RECT 1.780 2.115 1.950 2.285 ;
        RECT 2.140 2.115 2.310 2.285 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_4

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 5.440 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.603000 ;
    PORT
      LAYER li1 ;
        RECT 2.970 1.070 3.290 1.540 ;
    END
  END A
  PIN LOWLVPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 1.920 1.305 2.980 4.135 ;
      LAYER met1 ;
        RECT 1.360 2.280 2.370 2.315 ;
        RECT 0.070 2.140 6.170 2.280 ;
        RECT 1.360 2.085 2.370 2.140 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 2.555 5.250 5.555 5.335 ;
        RECT 0.015 4.465 0.445 5.250 ;
        RECT 2.555 4.465 6.225 5.250 ;
        RECT 2.555 4.425 5.555 4.465 ;
      LAYER met1 ;
        RECT 0.000 5.200 6.440 5.680 ;
    END
    PORT
      LAYER pwell ;
        RECT 3.005 0.975 5.705 1.070 ;
        RECT 0.015 0.190 0.445 0.975 ;
        RECT 3.005 0.960 6.225 0.975 ;
        RECT 1.990 0.280 6.225 0.960 ;
        RECT 3.005 0.190 6.225 0.280 ;
        RECT 3.005 0.160 5.705 0.190 ;
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 4.135 ;
        RECT 4.250 1.305 6.630 4.135 ;
      LAYER met1 ;
        RECT 0.080 3.640 0.370 3.685 ;
        RECT 5.870 3.640 6.160 3.685 ;
        RECT 0.070 3.500 6.170 3.640 ;
        RECT 0.080 3.455 0.370 3.500 ;
        RECT 5.870 3.455 6.160 3.500 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.402500 ;
    PORT
      LAYER li1 ;
        RECT 5.360 0.980 5.635 2.370 ;
        RECT 5.335 0.290 5.635 0.980 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 5.355 6.440 5.525 ;
        RECT 0.085 4.630 0.375 5.355 ;
        RECT 2.645 4.515 2.905 5.355 ;
        RECT 3.075 4.325 3.405 5.185 ;
        RECT 3.575 4.515 3.765 5.355 ;
        RECT 3.935 4.325 4.265 5.185 ;
        RECT 4.445 4.515 4.955 5.355 ;
        RECT 5.135 4.820 5.485 5.160 ;
        RECT 5.135 4.460 5.695 4.820 ;
        RECT 5.865 4.630 6.155 5.355 ;
        RECT 5.135 4.405 5.765 4.460 ;
        RECT 3.075 4.265 4.265 4.325 ;
        RECT 5.360 4.355 5.765 4.405 ;
        RECT 3.145 4.155 4.195 4.265 ;
        RECT 0.085 2.985 0.375 3.970 ;
        RECT 0.000 2.635 1.890 2.805 ;
        RECT 2.060 2.660 2.810 3.750 ;
        RECT 2.060 2.335 2.390 2.660 ;
        RECT 3.060 2.370 3.390 3.965 ;
        RECT 4.020 3.810 4.190 4.155 ;
        RECT 5.360 4.125 6.085 4.355 ;
        RECT 4.410 3.640 4.720 3.740 ;
        RECT 3.680 3.470 4.720 3.640 ;
        RECT 3.680 2.575 3.850 3.470 ;
        RECT 4.020 2.915 4.190 3.300 ;
        RECT 4.390 3.085 4.720 3.470 ;
        RECT 4.020 2.745 4.640 2.915 ;
        RECT 3.680 2.405 4.190 2.575 ;
        RECT 1.380 2.065 2.390 2.335 ;
        RECT 2.060 1.635 2.390 2.065 ;
        RECT 2.560 2.130 3.390 2.370 ;
        RECT 0.085 0.085 0.375 0.810 ;
        RECT 2.020 0.085 2.350 0.895 ;
        RECT 2.560 0.375 2.800 2.130 ;
        RECT 4.020 0.980 4.190 2.405 ;
        RECT 4.470 1.625 4.640 2.745 ;
        RECT 4.890 2.805 5.120 3.740 ;
        RECT 5.360 3.070 5.550 4.125 ;
        RECT 5.865 2.985 6.155 3.955 ;
        RECT 4.890 2.635 6.440 2.805 ;
        RECT 4.890 1.625 5.120 2.635 ;
        RECT 3.115 0.085 3.445 0.900 ;
        RECT 3.615 0.730 4.665 0.980 ;
        RECT 3.615 0.290 3.805 0.730 ;
        RECT 3.975 0.085 4.305 0.560 ;
        RECT 4.475 0.290 4.665 0.730 ;
        RECT 4.835 0.085 5.165 0.900 ;
        RECT 5.865 0.085 6.155 0.810 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 5.355 0.315 5.525 ;
        RECT 0.605 5.355 0.775 5.525 ;
        RECT 1.065 5.355 1.235 5.525 ;
        RECT 1.525 5.355 1.695 5.525 ;
        RECT 1.985 5.355 2.155 5.525 ;
        RECT 2.445 5.355 2.615 5.525 ;
        RECT 2.905 5.355 3.075 5.525 ;
        RECT 3.365 5.355 3.535 5.525 ;
        RECT 3.825 5.355 3.995 5.525 ;
        RECT 4.285 5.355 4.455 5.525 ;
        RECT 4.745 5.355 4.915 5.525 ;
        RECT 5.205 5.355 5.375 5.525 ;
        RECT 5.665 5.355 5.835 5.525 ;
        RECT 6.125 5.355 6.295 5.525 ;
        RECT 0.140 3.485 0.310 3.655 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.420 2.115 1.590 2.285 ;
        RECT 1.780 2.115 1.950 2.285 ;
        RECT 2.140 2.115 2.310 2.285 ;
        RECT 5.930 3.485 6.100 3.655 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_1

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 5.440 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.603000 ;
    PORT
      LAYER li1 ;
        RECT 2.970 1.070 3.290 1.540 ;
    END
  END A
  PIN LOWLVPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 1.920 1.305 2.980 4.135 ;
      LAYER met1 ;
        RECT 1.360 2.280 2.370 2.315 ;
        RECT 0.070 2.140 6.370 2.280 ;
        RECT 1.360 2.085 2.370 2.140 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 2.555 5.250 5.555 5.335 ;
        RECT 0.015 4.465 0.445 5.250 ;
        RECT 2.555 4.465 6.425 5.250 ;
        RECT 2.555 4.425 5.555 4.465 ;
      LAYER met1 ;
        RECT 0.000 5.200 6.440 5.680 ;
    END
    PORT
      LAYER pwell ;
        RECT 0.015 0.190 0.445 0.975 ;
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 4.135 ;
        RECT 4.250 1.305 6.630 4.135 ;
      LAYER met1 ;
        RECT 0.080 3.640 0.370 3.685 ;
        RECT 6.010 3.640 6.300 3.685 ;
        RECT 0.070 3.500 6.300 3.640 ;
        RECT 0.080 3.455 0.370 3.500 ;
        RECT 6.010 3.455 6.300 3.500 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.610500 ;
    PORT
      LAYER li1 ;
        RECT 5.360 0.980 5.635 2.370 ;
        RECT 5.335 0.255 5.635 0.980 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 3.005 0.960 6.265 1.015 ;
        RECT 1.990 0.280 6.265 0.960 ;
        RECT 3.005 0.105 6.265 0.280 ;
      LAYER li1 ;
        RECT 0.000 5.355 6.440 5.525 ;
        RECT 0.085 4.630 0.375 5.355 ;
        RECT 2.645 4.515 2.905 5.355 ;
        RECT 3.075 4.325 3.405 5.185 ;
        RECT 3.575 4.515 3.765 5.355 ;
        RECT 3.935 4.325 4.265 5.185 ;
        RECT 4.445 4.515 4.955 5.355 ;
        RECT 5.135 4.820 5.485 5.160 ;
        RECT 5.135 4.460 5.695 4.820 ;
        RECT 6.065 4.630 6.355 5.355 ;
        RECT 5.135 4.405 5.765 4.460 ;
        RECT 3.075 4.265 4.265 4.325 ;
        RECT 5.360 4.355 5.765 4.405 ;
        RECT 3.145 4.155 4.195 4.265 ;
        RECT 0.085 2.985 0.375 3.970 ;
        RECT 0.000 2.635 1.890 2.805 ;
        RECT 2.060 2.660 2.810 3.750 ;
        RECT 2.060 2.335 2.390 2.660 ;
        RECT 3.060 2.370 3.390 3.965 ;
        RECT 4.020 3.810 4.190 4.155 ;
        RECT 5.360 4.125 6.085 4.355 ;
        RECT 4.410 3.640 4.720 3.740 ;
        RECT 3.680 3.470 4.720 3.640 ;
        RECT 3.680 2.575 3.850 3.470 ;
        RECT 4.020 2.915 4.190 3.300 ;
        RECT 4.390 3.085 4.720 3.470 ;
        RECT 4.020 2.745 4.640 2.915 ;
        RECT 3.680 2.405 4.190 2.575 ;
        RECT 1.380 2.065 2.390 2.335 ;
        RECT 2.060 1.635 2.390 2.065 ;
        RECT 2.560 2.130 3.390 2.370 ;
        RECT 0.085 0.085 0.375 0.810 ;
        RECT 2.020 0.085 2.350 0.895 ;
        RECT 2.560 0.375 2.800 2.130 ;
        RECT 4.020 0.980 4.190 2.405 ;
        RECT 4.470 1.625 4.640 2.745 ;
        RECT 4.890 2.805 5.120 3.740 ;
        RECT 5.360 3.070 5.550 4.125 ;
        RECT 6.065 2.985 6.355 3.955 ;
        RECT 4.890 2.635 6.440 2.805 ;
        RECT 4.890 1.625 5.120 2.635 ;
        RECT 5.905 1.610 6.075 2.635 ;
        RECT 3.115 0.085 3.445 0.900 ;
        RECT 3.615 0.730 4.665 0.980 ;
        RECT 3.615 0.255 3.805 0.730 ;
        RECT 3.975 0.085 4.305 0.560 ;
        RECT 4.475 0.255 4.665 0.730 ;
        RECT 4.835 0.085 5.165 0.900 ;
        RECT 5.825 0.085 6.155 0.900 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 5.355 0.315 5.525 ;
        RECT 0.605 5.355 0.775 5.525 ;
        RECT 1.065 5.355 1.235 5.525 ;
        RECT 1.525 5.355 1.695 5.525 ;
        RECT 1.985 5.355 2.155 5.525 ;
        RECT 2.445 5.355 2.615 5.525 ;
        RECT 2.905 5.355 3.075 5.525 ;
        RECT 3.365 5.355 3.535 5.525 ;
        RECT 3.825 5.355 3.995 5.525 ;
        RECT 4.285 5.355 4.455 5.525 ;
        RECT 4.745 5.355 4.915 5.525 ;
        RECT 5.205 5.355 5.375 5.525 ;
        RECT 5.665 5.355 5.835 5.525 ;
        RECT 6.125 5.355 6.295 5.525 ;
        RECT 0.140 3.485 0.310 3.655 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.420 2.115 1.590 2.285 ;
        RECT 1.780 2.115 1.950 2.285 ;
        RECT 2.140 2.115 2.310 2.285 ;
        RECT 6.070 3.485 6.240 3.655 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_2

#--------EOF---------

MACRO sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 5.440 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.603000 ;
    PORT
      LAYER li1 ;
        RECT 2.970 1.070 3.290 1.540 ;
    END
  END A
  PIN LOWLVPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 1.920 1.305 2.980 4.135 ;
      LAYER met1 ;
        RECT 1.360 2.280 2.370 2.315 ;
        RECT 0.070 2.140 7.290 2.280 ;
        RECT 1.360 2.085 2.370 2.140 ;
    END
  END LOWLVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 0.015 4.465 0.445 5.250 ;
        RECT 6.915 4.465 7.345 5.250 ;
      LAYER met1 ;
        RECT 0.000 5.200 7.360 5.680 ;
    END
    PORT
      LAYER pwell ;
        RECT 0.015 0.190 0.445 0.975 ;
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 4.135 ;
        RECT 4.250 1.305 7.405 4.135 ;
      LAYER met1 ;
        RECT 0.080 3.640 0.370 3.685 ;
        RECT 6.930 3.640 7.220 3.685 ;
        RECT 0.070 3.500 7.290 3.640 ;
        RECT 0.080 3.455 0.370 3.500 ;
        RECT 6.930 3.455 7.220 3.500 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.072500 ;
    PORT
      LAYER li1 ;
        RECT 5.360 1.410 5.635 2.370 ;
        RECT 6.280 1.410 6.555 2.370 ;
        RECT 5.360 1.085 6.555 1.410 ;
        RECT 5.360 0.980 5.635 1.085 ;
        RECT 5.335 0.255 5.635 0.980 ;
        RECT 6.335 0.255 6.555 1.085 ;
    END
  END X
  OBS
      LAYER pwell ;
        RECT 2.555 4.425 5.555 5.335 ;
        RECT 3.005 0.960 7.125 1.015 ;
        RECT 1.990 0.280 7.125 0.960 ;
        RECT 3.005 0.105 7.125 0.280 ;
      LAYER li1 ;
        RECT 0.000 5.355 7.360 5.525 ;
        RECT 0.085 4.630 0.375 5.355 ;
        RECT 2.645 4.515 2.905 5.355 ;
        RECT 3.075 4.325 3.405 5.185 ;
        RECT 3.575 4.515 3.765 5.355 ;
        RECT 3.935 4.325 4.265 5.185 ;
        RECT 4.445 4.515 4.955 5.355 ;
        RECT 5.135 4.820 5.485 5.160 ;
        RECT 5.135 4.460 5.695 4.820 ;
        RECT 6.985 4.630 7.275 5.355 ;
        RECT 5.135 4.405 5.765 4.460 ;
        RECT 3.075 4.265 4.265 4.325 ;
        RECT 5.360 4.355 5.765 4.405 ;
        RECT 3.145 4.155 4.195 4.265 ;
        RECT 0.085 2.985 0.375 3.970 ;
        RECT 0.000 2.635 1.890 2.805 ;
        RECT 2.060 2.660 2.810 3.750 ;
        RECT 2.060 2.335 2.390 2.660 ;
        RECT 3.060 2.370 3.390 3.965 ;
        RECT 4.020 3.810 4.190 4.155 ;
        RECT 5.360 4.125 6.085 4.355 ;
        RECT 4.410 3.640 4.720 3.740 ;
        RECT 3.680 3.470 4.720 3.640 ;
        RECT 3.680 2.575 3.850 3.470 ;
        RECT 4.020 2.915 4.190 3.300 ;
        RECT 4.390 3.085 4.720 3.470 ;
        RECT 4.020 2.745 4.640 2.915 ;
        RECT 3.680 2.405 4.190 2.575 ;
        RECT 1.380 2.065 2.390 2.335 ;
        RECT 2.060 1.635 2.390 2.065 ;
        RECT 2.560 2.130 3.390 2.370 ;
        RECT 0.085 0.085 0.375 0.810 ;
        RECT 2.020 0.085 2.350 0.895 ;
        RECT 2.560 0.375 2.800 2.130 ;
        RECT 4.020 0.980 4.190 2.405 ;
        RECT 4.470 1.625 4.640 2.745 ;
        RECT 4.890 2.805 5.120 3.740 ;
        RECT 5.360 3.070 5.550 4.125 ;
        RECT 6.985 2.985 7.275 3.955 ;
        RECT 4.890 2.635 7.360 2.805 ;
        RECT 4.890 1.625 5.120 2.635 ;
        RECT 5.905 1.610 6.075 2.635 ;
        RECT 6.755 1.610 6.935 2.635 ;
        RECT 3.115 0.085 3.445 0.900 ;
        RECT 3.615 0.730 4.665 0.980 ;
        RECT 3.615 0.255 3.805 0.730 ;
        RECT 3.975 0.085 4.305 0.560 ;
        RECT 4.475 0.255 4.665 0.730 ;
        RECT 4.835 0.085 5.165 0.900 ;
        RECT 5.825 0.085 6.155 0.845 ;
        RECT 6.755 0.085 7.005 0.925 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 5.355 0.315 5.525 ;
        RECT 0.605 5.355 0.775 5.525 ;
        RECT 1.065 5.355 1.235 5.525 ;
        RECT 1.525 5.355 1.695 5.525 ;
        RECT 1.985 5.355 2.155 5.525 ;
        RECT 2.445 5.355 2.615 5.525 ;
        RECT 2.905 5.355 3.075 5.525 ;
        RECT 3.365 5.355 3.535 5.525 ;
        RECT 3.825 5.355 3.995 5.525 ;
        RECT 4.285 5.355 4.455 5.525 ;
        RECT 4.745 5.355 4.915 5.525 ;
        RECT 5.205 5.355 5.375 5.525 ;
        RECT 5.665 5.355 5.835 5.525 ;
        RECT 6.125 5.355 6.295 5.525 ;
        RECT 6.585 5.355 6.755 5.525 ;
        RECT 7.045 5.355 7.215 5.525 ;
        RECT 0.140 3.485 0.310 3.655 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.420 2.115 1.590 2.285 ;
        RECT 1.780 2.115 1.950 2.285 ;
        RECT 2.140 2.115 2.310 2.285 ;
        RECT 6.990 3.485 7.160 3.655 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
END sky130_fd_sc_hd__lpflow_lsbuf_lh_isowell_tap_4

#--------EOF---------

MACRO sky130_fd_sc_hd__macro_sparecell
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__macro_sparecell ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.340 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 13.340 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 13.530 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 13.340 2.960 ;
    END
  END VPWR
  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER met1 ;
        RECT 4.715 1.260 5.005 1.305 ;
        RECT 5.645 1.260 5.935 1.305 ;
        RECT 6.705 1.260 6.995 1.305 ;
        RECT 7.565 1.260 7.855 1.305 ;
        RECT 8.425 1.260 8.715 1.305 ;
        RECT 4.715 1.120 8.715 1.260 ;
        RECT 4.715 1.075 5.005 1.120 ;
        RECT 5.645 1.075 5.935 1.120 ;
        RECT 6.705 1.075 6.995 1.120 ;
        RECT 7.565 1.075 7.855 1.120 ;
        RECT 8.425 1.075 8.715 1.120 ;
    END
  END LO
  OBS
      LAYER pwell ;
        RECT 0.015 0.105 1.365 1.015 ;
        RECT 1.465 0.105 3.675 1.015 ;
        RECT 3.785 0.105 5.975 1.015 ;
        RECT 7.365 0.105 9.555 1.015 ;
        RECT 9.665 0.105 11.875 1.015 ;
        RECT 11.975 0.105 13.325 1.015 ;
        RECT 1.065 -0.085 1.235 0.105 ;
        RECT 3.360 -0.085 3.530 0.105 ;
        RECT 5.660 -0.085 5.830 0.105 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 7.510 -0.085 7.680 0.105 ;
        RECT 9.810 -0.085 9.980 0.105 ;
        RECT 12.105 -0.085 12.275 0.105 ;
      LAYER li1 ;
        RECT 0.000 2.635 13.340 2.805 ;
        RECT 0.145 1.495 0.355 2.635 ;
        RECT 0.525 1.485 0.855 2.465 ;
        RECT 1.025 1.495 1.255 2.635 ;
        RECT 1.505 2.295 2.645 2.465 ;
        RECT 1.505 1.835 1.805 2.295 ;
        RECT 1.975 1.665 2.305 2.125 ;
        RECT 0.145 0.085 0.355 0.905 ;
        RECT 0.525 0.885 0.775 1.485 ;
        RECT 1.545 1.445 2.305 1.665 ;
        RECT 2.475 1.665 2.645 2.295 ;
        RECT 2.815 1.835 3.145 2.635 ;
        RECT 3.315 1.665 3.590 2.465 ;
        RECT 3.870 1.835 4.125 2.635 ;
        RECT 4.295 1.665 4.625 2.465 ;
        RECT 4.795 1.835 4.965 2.635 ;
        RECT 5.135 1.665 5.465 2.465 ;
        RECT 2.475 1.455 3.590 1.665 ;
        RECT 3.765 1.495 5.465 1.665 ;
        RECT 5.635 1.495 5.895 2.635 ;
        RECT 6.255 1.910 6.585 2.635 ;
        RECT 0.945 1.075 1.275 1.325 ;
        RECT 1.545 0.905 1.760 1.445 ;
        RECT 1.930 1.075 2.700 1.275 ;
        RECT 2.870 1.075 3.590 1.275 ;
        RECT 3.765 0.905 4.045 1.495 ;
        RECT 4.215 1.075 4.965 1.325 ;
        RECT 5.135 1.075 5.895 1.325 ;
        RECT 0.525 0.255 0.855 0.885 ;
        RECT 1.025 0.085 1.255 0.905 ;
        RECT 1.545 0.735 3.145 0.905 ;
        RECT 1.975 0.725 3.145 0.735 ;
        RECT 1.515 0.085 1.805 0.555 ;
        RECT 1.975 0.255 2.305 0.725 ;
        RECT 2.475 0.085 2.645 0.555 ;
        RECT 2.815 0.255 3.145 0.725 ;
        RECT 3.315 0.085 3.590 0.905 ;
        RECT 3.765 0.655 4.625 0.905 ;
        RECT 4.795 0.715 5.895 0.885 ;
        RECT 3.875 0.465 4.205 0.485 ;
        RECT 4.795 0.465 5.045 0.715 ;
        RECT 3.875 0.255 5.045 0.465 ;
        RECT 5.215 0.085 5.385 0.545 ;
        RECT 5.555 0.255 5.895 0.715 ;
        RECT 6.065 0.255 6.585 1.740 ;
        RECT 6.755 0.915 7.275 2.465 ;
        RECT 7.445 1.495 7.705 2.635 ;
        RECT 7.875 1.665 8.205 2.465 ;
        RECT 8.375 1.835 8.545 2.635 ;
        RECT 8.715 1.665 9.045 2.465 ;
        RECT 9.215 1.835 9.470 2.635 ;
        RECT 9.750 1.665 10.025 2.465 ;
        RECT 10.195 1.835 10.525 2.635 ;
        RECT 10.695 2.295 11.835 2.465 ;
        RECT 10.695 1.665 10.865 2.295 ;
        RECT 7.875 1.495 9.575 1.665 ;
        RECT 7.445 1.075 8.205 1.325 ;
        RECT 8.375 1.075 9.125 1.325 ;
        RECT 9.295 0.905 9.575 1.495 ;
        RECT 9.750 1.455 10.865 1.665 ;
        RECT 11.035 1.665 11.365 2.125 ;
        RECT 11.535 1.835 11.835 2.295 ;
        RECT 11.035 1.445 11.795 1.665 ;
        RECT 12.085 1.495 12.315 2.635 ;
        RECT 12.485 1.485 12.815 2.465 ;
        RECT 12.985 1.495 13.195 2.635 ;
        RECT 9.750 1.075 10.470 1.275 ;
        RECT 10.640 1.075 11.410 1.275 ;
        RECT 11.580 0.905 11.795 1.445 ;
        RECT 12.065 1.075 12.395 1.325 ;
        RECT 6.755 0.085 7.095 0.745 ;
        RECT 7.445 0.715 8.545 0.885 ;
        RECT 7.445 0.255 7.785 0.715 ;
        RECT 7.955 0.085 8.125 0.545 ;
        RECT 8.295 0.465 8.545 0.715 ;
        RECT 8.715 0.655 9.575 0.905 ;
        RECT 9.135 0.465 9.465 0.485 ;
        RECT 8.295 0.255 9.465 0.465 ;
        RECT 9.750 0.085 10.025 0.905 ;
        RECT 10.195 0.735 11.795 0.905 ;
        RECT 10.195 0.725 11.365 0.735 ;
        RECT 10.195 0.255 10.525 0.725 ;
        RECT 10.695 0.085 10.865 0.555 ;
        RECT 11.035 0.255 11.365 0.725 ;
        RECT 11.535 0.085 11.825 0.555 ;
        RECT 12.085 0.085 12.315 0.905 ;
        RECT 12.565 0.885 12.815 1.485 ;
        RECT 12.485 0.255 12.815 0.885 ;
        RECT 12.985 0.085 13.195 0.905 ;
        RECT 0.000 -0.085 13.340 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 0.565 1.105 0.735 1.275 ;
        RECT 1.085 1.105 1.255 1.275 ;
        RECT 1.570 1.105 1.740 1.275 ;
        RECT 2.100 1.105 2.270 1.275 ;
        RECT 2.960 1.105 3.130 1.275 ;
        RECT 3.820 1.105 3.990 1.275 ;
        RECT 4.775 1.105 4.945 1.275 ;
        RECT 5.705 1.105 5.875 1.275 ;
        RECT 6.765 1.105 6.935 1.275 ;
        RECT 7.625 1.105 7.795 1.275 ;
        RECT 8.485 1.105 8.655 1.275 ;
        RECT 9.345 1.105 9.515 1.275 ;
        RECT 10.205 1.105 10.375 1.275 ;
        RECT 11.065 1.105 11.235 1.275 ;
        RECT 11.605 1.105 11.775 1.275 ;
        RECT 12.090 1.105 12.260 1.275 ;
        RECT 12.605 1.105 12.775 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
      LAYER met1 ;
        RECT 0.505 1.075 0.875 1.305 ;
        RECT 1.025 1.260 1.315 1.305 ;
        RECT 1.510 1.260 1.800 1.305 ;
        RECT 1.025 1.120 1.800 1.260 ;
        RECT 1.025 1.075 1.315 1.120 ;
        RECT 1.510 1.075 1.800 1.120 ;
        RECT 2.040 1.260 2.330 1.305 ;
        RECT 2.900 1.260 3.190 1.305 ;
        RECT 3.760 1.260 4.050 1.305 ;
        RECT 2.040 1.120 4.050 1.260 ;
        RECT 2.040 1.075 2.330 1.120 ;
        RECT 2.900 1.075 3.190 1.120 ;
        RECT 3.760 1.075 4.050 1.120 ;
        RECT 9.285 1.260 9.575 1.305 ;
        RECT 10.145 1.260 10.435 1.305 ;
        RECT 11.005 1.260 11.295 1.305 ;
        RECT 9.285 1.120 11.295 1.260 ;
        RECT 9.285 1.075 9.575 1.120 ;
        RECT 10.145 1.075 10.435 1.120 ;
        RECT 11.005 1.075 11.295 1.120 ;
        RECT 11.545 1.260 11.835 1.305 ;
        RECT 12.030 1.260 12.320 1.305 ;
        RECT 11.545 1.120 12.320 1.260 ;
        RECT 11.545 1.075 11.835 1.120 ;
        RECT 12.030 1.075 12.320 1.120 ;
        RECT 12.470 1.075 12.835 1.305 ;
  END
END sky130_fd_sc_hd__macro_sparecell

#--------EOF---------

MACRO sky130_fd_sc_hd__maj3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__maj3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT 0.610 1.325 0.780 2.460 ;
        RECT 0.610 0.995 1.125 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT 1.500 0.995 1.905 1.615 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT 2.415 0.765 2.755 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.650 0.785 3.675 1.015 ;
        RECT 0.005 0.105 3.675 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.602250 ;
    PORT
      LAYER li1 ;
        RECT 3.255 2.160 3.595 2.465 ;
        RECT 3.265 1.495 3.595 2.160 ;
        RECT 3.370 0.825 3.595 1.495 ;
        RECT 3.255 0.255 3.595 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.135 0.825 0.395 2.125 ;
        RECT 0.955 1.715 1.205 2.635 ;
        RECT 1.655 1.815 2.245 2.080 ;
        RECT 2.555 1.845 2.885 2.635 ;
        RECT 2.075 1.665 2.245 1.815 ;
        RECT 2.075 1.495 3.095 1.665 ;
        RECT 2.075 0.825 2.245 1.495 ;
        RECT 2.925 1.325 3.095 1.495 ;
        RECT 2.925 0.995 3.200 1.325 ;
        RECT 0.135 0.655 2.245 0.825 ;
        RECT 0.135 0.255 0.395 0.655 ;
        RECT 1.655 0.640 2.245 0.655 ;
        RECT 0.875 0.085 1.205 0.485 ;
        RECT 1.655 0.255 1.985 0.640 ;
        RECT 2.545 0.085 2.880 0.470 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__maj3_1

#--------EOF---------

MACRO sky130_fd_sc_hd__maj3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__maj3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 1.005 0.995 1.695 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 1.865 0.995 2.155 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.495 3.070 1.665 ;
        RECT 0.425 0.995 0.775 1.495 ;
        RECT 2.415 1.415 3.070 1.495 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.720 0.785 4.135 1.015 ;
        RECT 0.105 0.105 4.135 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 3.285 1.495 3.615 2.465 ;
        RECT 3.445 0.905 3.615 1.495 ;
        RECT 3.285 0.255 3.615 0.905 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 2.005 0.615 2.465 ;
        RECT 0.975 2.175 1.305 2.635 ;
        RECT 1.755 2.005 2.085 2.465 ;
        RECT 0.085 1.835 2.085 2.005 ;
        RECT 2.535 1.835 2.860 2.635 ;
        RECT 0.085 0.825 0.255 1.835 ;
        RECT 3.785 1.495 4.055 2.635 ;
        RECT 2.925 1.075 3.275 1.245 ;
        RECT 2.925 0.825 3.105 1.075 ;
        RECT 0.085 0.655 3.105 0.825 ;
        RECT 0.085 0.280 0.525 0.655 ;
        RECT 0.975 0.085 1.305 0.485 ;
        RECT 1.755 0.255 2.085 0.655 ;
        RECT 2.635 0.085 2.965 0.485 ;
        RECT 3.785 0.085 4.055 0.905 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__maj3_2

#--------EOF---------

MACRO sky130_fd_sc_hd__maj3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__maj3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.060 1.075 1.450 1.635 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.960 1.075 2.290 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.620 2.225 2.630 2.395 ;
        RECT 1.620 2.085 1.790 2.225 ;
        RECT 0.720 1.915 1.790 2.085 ;
        RECT 0.720 1.285 0.890 1.915 ;
        RECT 0.425 1.075 0.890 1.285 ;
        RECT 2.460 1.245 2.630 2.225 ;
        RECT 2.460 1.075 2.945 1.245 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.195 0.105 5.055 1.015 ;
        RECT 0.195 0.085 0.310 0.105 ;
        RECT 0.140 -0.085 0.310 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 3.375 1.625 3.705 2.465 ;
        RECT 4.215 1.625 4.545 2.465 ;
        RECT 3.375 1.455 4.975 1.625 ;
        RECT 4.715 0.905 4.975 1.455 ;
        RECT 3.455 0.715 4.975 0.905 ;
        RECT 3.455 0.490 3.705 0.715 ;
        RECT 3.375 0.255 3.705 0.490 ;
        RECT 4.215 0.255 4.545 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.085 1.455 0.465 2.465 ;
        RECT 1.120 2.255 1.450 2.635 ;
        RECT 1.960 1.745 2.290 2.055 ;
        RECT 1.620 1.545 2.290 1.745 ;
        RECT 0.085 0.885 0.255 1.455 ;
        RECT 1.620 0.885 1.790 1.545 ;
        RECT 2.845 1.455 3.175 2.635 ;
        RECT 3.875 1.795 4.045 2.635 ;
        RECT 4.715 1.795 4.925 2.635 ;
        RECT 3.115 1.075 4.545 1.285 ;
        RECT 3.115 0.885 3.285 1.075 ;
        RECT 0.085 0.715 3.285 0.885 ;
        RECT 0.085 0.660 2.290 0.715 ;
        RECT 0.085 0.255 0.635 0.660 ;
        RECT 1.120 0.085 1.450 0.490 ;
        RECT 1.960 0.255 2.290 0.660 ;
        RECT 2.860 0.085 3.205 0.545 ;
        RECT 3.875 0.085 4.045 0.545 ;
        RECT 4.715 0.085 4.885 0.545 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
END sky130_fd_sc_hd__maj3_4

#--------EOF---------

MACRO sky130_fd_sc_hd__mux2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.990 0.255 2.265 1.415 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.615 1.615 2.625 1.785 ;
        RECT 1.615 0.815 1.785 1.615 ;
        RECT 2.435 0.255 2.625 1.615 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT 0.935 2.295 2.965 2.465 ;
        RECT 0.935 1.325 1.105 2.295 ;
        RECT 2.795 1.630 2.965 2.295 ;
        RECT 2.795 1.440 3.545 1.630 ;
        RECT 0.910 0.995 1.105 1.325 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 0.935 1.015 ;
        RECT 0.005 0.105 3.905 0.785 ;
        RECT 0.420 -0.085 0.590 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.495 0.425 2.465 ;
        RECT 0.090 0.825 0.260 1.495 ;
        RECT 0.090 0.255 0.345 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.595 1.495 0.765 2.635 ;
        RECT 1.275 1.955 2.400 2.125 ;
        RECT 0.430 0.995 0.685 1.325 ;
        RECT 0.515 0.825 0.685 0.995 ;
        RECT 1.275 0.825 1.445 1.955 ;
        RECT 3.135 1.875 3.305 2.635 ;
        RECT 3.540 1.875 4.055 2.285 ;
        RECT 3.715 1.065 4.055 1.875 ;
        RECT 2.825 0.895 4.055 1.065 ;
        RECT 0.515 0.655 1.445 0.825 ;
        RECT 1.270 0.620 1.445 0.655 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.270 0.255 1.800 0.620 ;
        RECT 2.805 0.085 3.315 0.620 ;
        RECT 3.535 0.290 3.780 0.895 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__mux2_1

#--------EOF---------

MACRO sky130_fd_sc_hd__mux2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.275 1.315 3.090 1.625 ;
        RECT 2.275 1.280 2.445 1.315 ;
        RECT 1.815 0.765 2.445 1.280 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.625 0.735 3.090 1.025 ;
        RECT 2.900 0.420 3.090 0.735 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 3.360 0.755 3.550 1.625 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 1.345 1.015 ;
        RECT 0.005 0.105 4.135 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.595 0.825 2.465 ;
        RECT 0.515 0.750 0.685 1.595 ;
        RECT 0.515 0.255 0.765 0.750 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.025 2.175 1.315 2.635 ;
        RECT 1.485 2.255 2.795 2.425 ;
        RECT 1.485 2.005 1.655 2.255 ;
        RECT 3.325 2.175 3.545 2.635 ;
        RECT 3.715 2.005 4.050 2.465 ;
        RECT 0.995 1.835 1.655 2.005 ;
        RECT 1.825 1.835 4.050 2.005 ;
        RECT 0.995 1.325 1.165 1.835 ;
        RECT 1.825 1.665 1.995 1.835 ;
        RECT 0.855 0.995 1.165 1.325 ;
        RECT 1.335 1.495 1.995 1.665 ;
        RECT 1.335 0.995 1.505 1.495 ;
        RECT 0.090 0.085 0.345 0.885 ;
        RECT 0.995 0.805 1.165 0.995 ;
        RECT 0.995 0.635 1.605 0.805 ;
        RECT 1.435 0.465 1.605 0.635 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 1.435 0.295 2.730 0.465 ;
        RECT 3.350 0.085 3.550 0.585 ;
        RECT 3.720 0.255 4.050 1.835 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__mux2_2

#--------EOF---------

MACRO sky130_fd_sc_hd__mux2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.480 0.995 1.750 1.615 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.965 0.995 2.435 1.325 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.430 0.995 0.740 1.325 ;
        RECT 0.570 0.805 0.740 0.995 ;
        RECT 2.680 0.995 3.395 1.325 ;
        RECT 2.680 0.805 2.850 0.995 ;
        RECT 0.570 0.635 2.850 0.805 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.515 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 3.915 1.745 4.085 2.465 ;
        RECT 4.755 1.745 4.925 2.465 ;
        RECT 3.915 1.575 5.430 1.745 ;
        RECT 5.200 0.805 5.430 1.575 ;
        RECT 3.915 0.635 5.430 0.805 ;
        RECT 3.915 0.255 4.085 0.635 ;
        RECT 4.755 0.255 4.925 0.635 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.090 1.665 0.345 2.465 ;
        RECT 0.515 1.835 0.820 2.635 ;
        RECT 0.990 2.275 2.770 2.445 ;
        RECT 0.990 1.935 1.340 2.275 ;
        RECT 3.075 2.105 3.245 2.465 ;
        RECT 3.415 2.255 3.745 2.635 ;
        RECT 1.530 1.935 3.245 2.105 ;
        RECT 4.255 1.915 4.585 2.635 ;
        RECT 5.095 1.915 5.425 2.635 ;
        RECT 3.565 1.765 3.735 1.785 ;
        RECT 0.090 1.495 1.080 1.665 ;
        RECT 1.980 1.595 3.735 1.765 ;
        RECT 0.090 0.625 0.260 1.495 ;
        RECT 0.910 0.995 1.080 1.495 ;
        RECT 3.565 1.245 3.735 1.595 ;
        RECT 3.565 1.075 5.030 1.245 ;
        RECT 3.565 0.825 3.735 1.075 ;
        RECT 3.060 0.655 3.735 0.825 ;
        RECT 0.090 0.295 0.345 0.625 ;
        RECT 3.060 0.465 3.230 0.655 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.975 0.295 3.230 0.465 ;
        RECT 3.415 0.085 3.745 0.465 ;
        RECT 4.255 0.085 4.585 0.465 ;
        RECT 5.095 0.085 5.425 0.465 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__mux2_4

#--------EOF---------

MACRO sky130_fd_sc_hd__mux2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER li1 ;
        RECT 5.180 0.815 5.350 1.325 ;
        RECT 7.025 1.165 7.195 1.325 ;
        RECT 6.725 0.995 7.195 1.165 ;
        RECT 6.725 0.815 6.895 0.995 ;
        RECT 5.180 0.645 6.895 0.815 ;
        RECT 5.305 0.425 5.890 0.645 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492000 ;
    PORT
      LAYER met1 ;
        RECT 4.230 1.260 4.520 1.305 ;
        RECT 7.900 1.260 8.190 1.305 ;
        RECT 4.230 1.120 8.190 1.260 ;
        RECT 4.230 1.075 4.520 1.120 ;
        RECT 7.900 1.075 8.190 1.120 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.739500 ;
    PORT
      LAYER met1 ;
        RECT 5.610 1.600 5.900 1.645 ;
        RECT 9.280 1.600 9.570 1.645 ;
        RECT 5.610 1.460 9.570 1.600 ;
        RECT 5.610 1.415 5.900 1.460 ;
        RECT 9.280 1.415 9.570 1.460 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.005 3.865 1.015 ;
        RECT 8.735 1.005 9.655 1.015 ;
        RECT 0.005 0.105 9.655 1.005 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.745 0.765 2.465 ;
        RECT 1.435 1.745 1.605 2.465 ;
        RECT 2.275 1.745 2.445 2.465 ;
        RECT 3.115 1.745 3.285 2.465 ;
        RECT 0.595 1.575 3.285 1.745 ;
        RECT 0.595 0.805 0.815 1.575 ;
        RECT 0.595 0.635 3.285 0.805 ;
        RECT 0.595 0.255 0.765 0.635 ;
        RECT 1.435 0.295 1.605 0.635 ;
        RECT 2.275 0.255 2.445 0.635 ;
        RECT 3.115 0.295 3.285 0.635 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.090 1.915 0.425 2.635 ;
        RECT 0.935 1.915 1.265 2.635 ;
        RECT 1.775 1.915 2.105 2.635 ;
        RECT 2.615 1.915 2.945 2.635 ;
        RECT 3.455 2.255 3.785 2.635 ;
        RECT 3.955 2.255 5.905 2.425 ;
        RECT 6.075 2.175 6.245 2.635 ;
        RECT 6.480 2.255 8.645 2.425 ;
        RECT 8.815 2.255 9.145 2.635 ;
        RECT 9.315 2.085 9.485 2.465 ;
        RECT 3.455 1.835 8.225 2.005 ;
        RECT 8.685 1.915 9.485 2.085 ;
        RECT 3.455 1.245 3.625 1.835 ;
        RECT 8.685 1.665 8.855 1.915 ;
        RECT 9.315 1.795 9.485 1.915 ;
        RECT 0.985 1.075 3.625 1.245 ;
        RECT 3.455 0.805 3.625 1.075 ;
        RECT 3.795 1.495 6.035 1.665 ;
        RECT 3.795 0.995 3.965 1.495 ;
        RECT 4.305 1.275 4.475 1.325 ;
        RECT 4.290 1.105 4.475 1.275 ;
        RECT 4.305 0.995 4.475 1.105 ;
        RECT 5.670 0.995 6.035 1.495 ;
        RECT 6.345 1.495 8.855 1.665 ;
        RECT 6.345 0.995 6.515 1.495 ;
        RECT 7.960 0.995 8.245 1.325 ;
        RECT 4.750 0.805 4.920 0.935 ;
        RECT 7.500 0.805 7.670 0.935 ;
        RECT 3.455 0.635 4.920 0.805 ;
        RECT 7.115 0.635 7.670 0.805 ;
        RECT 8.685 0.815 8.855 1.495 ;
        RECT 9.215 0.995 9.510 1.615 ;
        RECT 8.685 0.645 9.485 0.815 ;
        RECT 0.090 0.085 0.425 0.465 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 1.775 0.085 2.105 0.465 ;
        RECT 2.615 0.085 2.945 0.465 ;
        RECT 3.455 0.085 3.785 0.465 ;
        RECT 3.955 0.295 5.125 0.465 ;
        RECT 6.060 0.085 6.390 0.465 ;
        RECT 6.575 0.295 7.865 0.465 ;
        RECT 8.815 0.085 9.145 0.465 ;
        RECT 9.315 0.295 9.485 0.645 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 5.670 1.445 5.840 1.615 ;
        RECT 4.290 1.105 4.460 1.275 ;
        RECT 7.960 1.105 8.130 1.275 ;
        RECT 4.750 0.765 4.920 0.935 ;
        RECT 7.500 0.765 7.670 0.935 ;
        RECT 9.340 1.445 9.510 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 4.690 0.920 4.980 0.965 ;
        RECT 7.440 0.920 7.730 0.965 ;
        RECT 4.690 0.780 7.730 0.920 ;
        RECT 4.690 0.735 4.980 0.780 ;
        RECT 7.440 0.735 7.730 0.780 ;
  END
END sky130_fd_sc_hd__mux2_8

#--------EOF---------

MACRO sky130_fd_sc_hd__mux2i_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2i_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.060 0.420 1.285 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.035 1.445 1.235 2.110 ;
        RECT 1.035 1.325 1.205 1.445 ;
        RECT 0.955 1.155 1.205 1.325 ;
        RECT 0.955 0.995 1.125 1.155 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.260 0.760 3.595 1.620 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.675 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.480500 ;
    PORT
      LAYER li1 ;
        RECT 0.590 1.455 0.840 2.125 ;
        RECT 0.590 0.595 0.780 1.455 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.120 2.295 1.575 2.465 ;
        RECT 0.120 1.455 0.420 2.295 ;
        RECT 1.405 1.650 1.575 2.295 ;
        RECT 1.745 1.835 1.975 2.635 ;
        RECT 2.285 1.650 2.615 2.465 ;
        RECT 1.405 1.480 2.615 1.650 ;
        RECT 2.860 1.310 3.085 2.465 ;
        RECT 3.295 1.835 3.590 2.635 ;
        RECT 1.385 1.075 3.085 1.310 ;
        RECT 0.085 0.465 0.345 0.885 ;
        RECT 1.295 0.825 2.620 0.885 ;
        RECT 0.955 0.715 2.620 0.825 ;
        RECT 0.955 0.655 1.520 0.715 ;
        RECT 0.085 0.425 0.440 0.465 ;
        RECT 0.965 0.425 1.805 0.465 ;
        RECT 0.085 0.255 1.805 0.425 ;
        RECT 1.975 0.085 2.145 0.545 ;
        RECT 2.385 0.255 2.620 0.715 ;
        RECT 2.800 0.485 3.085 1.075 ;
        RECT 2.800 0.255 3.165 0.485 ;
        RECT 3.335 0.085 3.555 0.545 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__mux2i_1

#--------EOF---------

MACRO sky130_fd_sc_hd__mux2i_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2i_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.470 1.075 3.560 1.275 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.310 0.995 4.635 1.615 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER li1 ;
        RECT 0.430 0.995 0.780 1.325 ;
        RECT 0.580 0.725 0.780 0.995 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.055 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.691250 ;
    PORT
      LAYER li1 ;
        RECT 2.715 2.255 4.975 2.425 ;
        RECT 4.750 1.785 4.975 2.255 ;
        RECT 4.805 0.465 4.975 1.785 ;
        RECT 2.715 0.295 4.975 0.465 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.085 2.135 0.345 2.465 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.355 2.255 1.685 2.635 ;
        RECT 1.855 2.135 2.080 2.465 ;
        RECT 2.275 2.175 2.525 2.635 ;
        RECT 0.085 1.665 0.260 2.135 ;
        RECT 1.910 2.005 2.080 2.135 ;
        RECT 2.715 2.005 4.350 2.085 ;
        RECT 0.935 1.835 1.735 2.005 ;
        RECT 1.910 1.915 4.350 2.005 ;
        RECT 1.910 1.835 2.885 1.915 ;
        RECT 1.565 1.665 1.735 1.835 ;
        RECT 3.135 1.665 3.465 1.715 ;
        RECT 0.085 1.495 1.395 1.665 ;
        RECT 1.565 1.495 3.465 1.665 ;
        RECT 0.085 0.675 0.260 1.495 ;
        RECT 1.225 1.325 1.395 1.495 ;
        RECT 1.225 1.155 1.985 1.325 ;
        RECT 1.655 1.075 1.985 1.155 ;
        RECT 0.085 0.345 0.345 0.675 ;
        RECT 1.015 0.575 1.255 0.935 ;
        RECT 0.515 0.085 0.835 0.545 ;
        RECT 1.435 0.085 1.685 0.885 ;
        RECT 1.855 0.735 3.465 0.905 ;
        RECT 1.855 0.295 2.025 0.735 ;
        RECT 3.135 0.655 3.465 0.735 ;
        RECT 3.850 0.825 4.105 0.935 ;
        RECT 3.850 0.655 4.345 0.825 ;
        RECT 2.275 0.085 2.445 0.545 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 1.070 0.765 1.240 0.935 ;
        RECT 3.850 0.765 4.020 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
      LAYER met1 ;
        RECT 1.010 0.920 1.300 0.965 ;
        RECT 3.790 0.920 4.080 0.965 ;
        RECT 1.010 0.780 4.080 0.920 ;
        RECT 1.010 0.735 1.300 0.780 ;
        RECT 3.790 0.735 4.080 0.780 ;
  END
END sky130_fd_sc_hd__mux2i_2

#--------EOF---------

MACRO sky130_fd_sc_hd__mux2i_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux2i_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.560 1.105 1.240 1.325 ;
        RECT 0.560 0.995 1.070 1.105 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.955 0.995 3.550 1.325 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.237500 ;
    PORT
      LAYER li1 ;
        RECT 5.760 1.425 7.850 1.595 ;
        RECT 5.760 1.290 5.930 1.425 ;
        RECT 3.845 1.075 5.930 1.290 ;
        RECT 7.680 0.995 7.850 1.425 ;
    END
  END S
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.275 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.194500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 2.255 3.785 2.425 ;
        RECT 0.095 0.485 0.320 2.255 ;
        RECT 0.095 0.315 3.785 0.485 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 3.975 2.255 4.305 2.635 ;
        RECT 4.815 2.255 5.145 2.635 ;
        RECT 5.655 2.255 5.985 2.635 ;
        RECT 6.155 2.085 6.325 2.465 ;
        RECT 6.495 2.255 6.825 2.635 ;
        RECT 6.995 2.085 7.165 2.465 ;
        RECT 7.435 2.255 7.765 2.635 ;
        RECT 2.195 1.915 7.165 2.085 ;
        RECT 6.155 1.795 6.325 1.915 ;
        RECT 6.995 1.795 7.165 1.915 ;
        RECT 7.935 1.795 8.195 2.465 ;
        RECT 0.515 1.575 5.580 1.745 ;
        RECT 6.730 1.075 7.510 1.245 ;
        RECT 1.355 0.825 1.700 0.935 ;
        RECT 6.150 0.905 6.450 0.935 ;
        RECT 0.515 0.655 1.700 0.825 ;
        RECT 2.195 0.655 5.485 0.825 ;
        RECT 3.975 0.085 4.305 0.465 ;
        RECT 4.475 0.255 4.645 0.655 ;
        RECT 4.815 0.085 5.145 0.465 ;
        RECT 5.315 0.255 5.485 0.655 ;
        RECT 6.150 0.715 7.165 0.905 ;
        RECT 5.655 0.085 5.980 0.590 ;
        RECT 6.150 0.255 6.325 0.715 ;
        RECT 6.545 0.085 6.795 0.545 ;
        RECT 6.995 0.510 7.165 0.715 ;
        RECT 7.340 0.825 7.510 1.075 ;
        RECT 8.020 0.825 8.195 1.795 ;
        RECT 7.340 0.655 8.195 0.825 ;
        RECT 7.435 0.085 7.765 0.465 ;
        RECT 7.935 0.255 8.195 0.655 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 1.530 0.765 1.700 0.935 ;
        RECT 6.150 0.765 6.320 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
      LAYER met1 ;
        RECT 1.470 0.920 1.760 0.965 ;
        RECT 6.090 0.920 6.380 0.965 ;
        RECT 1.470 0.780 6.380 0.920 ;
        RECT 1.470 0.735 1.760 0.780 ;
        RECT 6.090 0.735 6.380 0.780 ;
  END
END sky130_fd_sc_hd__mux2i_4

#--------EOF---------

MACRO sky130_fd_sc_hd__mux4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.805 0.995 1.240 1.615 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.150 0.995 0.495 1.615 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 5.250 1.055 5.580 1.675 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 4.800 1.055 5.045 1.675 ;
    END
  END A3
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER li1 ;
        RECT 3.265 0.995 3.565 1.995 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT 6.055 0.995 6.345 1.675 ;
    END
  END S1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 3.210 1.000 4.560 1.035 ;
        RECT 2.270 0.955 4.560 1.000 ;
        RECT 1.330 0.785 4.560 0.955 ;
        RECT 7.635 1.015 8.555 1.035 ;
        RECT 7.635 0.785 9.655 1.015 ;
        RECT 0.005 0.355 9.655 0.785 ;
        RECT 0.005 0.320 3.200 0.355 ;
        RECT 0.005 0.275 2.260 0.320 ;
        RECT 0.005 0.105 1.765 0.275 ;
        RECT 4.560 0.105 9.655 0.355 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 9.315 0.255 9.575 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.015 2.295 2.545 2.465 ;
        RECT 1.015 2.135 1.185 2.295 ;
        RECT 1.535 1.965 1.705 2.125 ;
        RECT 0.175 1.795 1.705 1.965 ;
        RECT 1.875 1.955 2.205 2.125 ;
        RECT 1.875 1.625 2.045 1.955 ;
        RECT 2.375 1.795 2.545 2.295 ;
        RECT 2.715 1.625 3.065 2.465 ;
        RECT 3.235 2.255 3.565 2.635 ;
        RECT 3.825 2.295 4.835 2.465 ;
        RECT 3.825 1.785 3.995 2.295 ;
        RECT 1.410 1.455 2.045 1.625 ;
        RECT 1.410 0.935 1.580 1.455 ;
        RECT 2.260 1.395 3.065 1.625 ;
        RECT 4.165 1.615 4.495 2.125 ;
        RECT 4.665 2.085 4.835 2.295 ;
        RECT 5.060 2.255 5.390 2.635 ;
        RECT 5.560 2.085 5.730 2.465 ;
        RECT 5.980 2.255 6.330 2.635 ;
        RECT 6.500 2.135 6.685 2.465 ;
        RECT 4.665 1.915 5.730 2.085 ;
        RECT 3.735 1.445 4.495 1.615 ;
        RECT 2.260 1.285 2.620 1.395 ;
        RECT 2.080 1.105 2.620 1.285 ;
        RECT 0.175 0.635 1.185 0.805 ;
        RECT 0.175 0.260 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.425 1.185 0.635 ;
        RECT 1.410 0.765 1.700 0.935 ;
        RECT 1.410 0.595 1.750 0.765 ;
        RECT 1.920 0.425 2.090 0.760 ;
        RECT 2.260 0.430 2.620 1.105 ;
        RECT 3.735 0.920 3.905 1.445 ;
        RECT 6.515 1.275 6.685 2.135 ;
        RECT 6.980 2.135 7.190 2.465 ;
        RECT 7.360 2.295 8.645 2.465 ;
        RECT 7.360 2.255 7.690 2.295 ;
        RECT 4.290 1.265 4.460 1.275 ;
        RECT 4.075 1.105 4.460 1.265 ;
        RECT 6.515 1.105 6.805 1.275 ;
        RECT 4.075 1.095 4.405 1.105 ;
        RECT 3.735 0.845 4.050 0.920 ;
        RECT 1.015 0.255 2.090 0.425 ;
        RECT 2.800 0.085 3.090 0.805 ;
        RECT 3.380 0.425 3.550 0.795 ;
        RECT 3.720 0.595 4.050 0.845 ;
        RECT 4.220 0.885 4.390 0.925 ;
        RECT 4.220 0.715 5.740 0.885 ;
        RECT 4.220 0.595 4.390 0.715 ;
        RECT 4.625 0.425 4.980 0.465 ;
        RECT 3.380 0.255 4.980 0.425 ;
        RECT 5.150 0.085 5.320 0.545 ;
        RECT 5.495 0.295 5.740 0.715 ;
        RECT 6.515 0.655 6.685 1.105 ;
        RECT 6.980 0.935 7.150 2.135 ;
        RECT 7.845 1.985 8.175 2.125 ;
        RECT 7.390 1.755 8.175 1.985 ;
        RECT 8.475 1.835 8.645 2.295 ;
        RECT 8.815 2.255 9.145 2.635 ;
        RECT 6.980 0.765 7.220 0.935 ;
        RECT 6.010 0.085 6.340 0.465 ;
        RECT 6.510 0.325 6.685 0.655 ;
        RECT 7.390 0.585 7.560 1.755 ;
        RECT 8.475 1.665 9.125 1.835 ;
        RECT 8.190 1.105 8.645 1.275 ;
        RECT 7.970 0.925 8.380 0.935 ;
        RECT 7.970 0.765 8.385 0.925 ;
        RECT 8.955 0.885 9.125 1.665 ;
        RECT 8.210 0.595 8.385 0.765 ;
        RECT 8.555 0.715 9.125 0.885 ;
        RECT 7.030 0.415 7.560 0.585 ;
        RECT 7.730 0.425 7.900 0.585 ;
        RECT 8.555 0.425 8.725 0.715 ;
        RECT 7.030 0.255 7.200 0.415 ;
        RECT 7.730 0.255 8.725 0.425 ;
        RECT 8.895 0.085 9.065 0.545 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 4.325 1.785 4.495 1.955 ;
        RECT 2.450 1.105 2.620 1.275 ;
        RECT 1.530 0.765 1.700 0.935 ;
        RECT 4.290 1.105 4.460 1.275 ;
        RECT 6.635 1.105 6.805 1.275 ;
        RECT 7.555 1.785 7.725 1.955 ;
        RECT 7.050 0.765 7.220 0.935 ;
        RECT 8.475 1.105 8.645 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 4.265 1.940 4.555 1.985 ;
        RECT 7.495 1.940 7.785 1.985 ;
        RECT 4.265 1.800 7.785 1.940 ;
        RECT 4.265 1.755 4.555 1.800 ;
        RECT 7.495 1.755 7.785 1.800 ;
        RECT 2.390 1.260 2.680 1.305 ;
        RECT 4.230 1.260 4.520 1.305 ;
        RECT 2.390 1.120 4.520 1.260 ;
        RECT 2.390 1.075 2.680 1.120 ;
        RECT 4.230 1.075 4.520 1.120 ;
        RECT 6.575 1.260 6.865 1.305 ;
        RECT 8.415 1.260 8.705 1.305 ;
        RECT 6.575 1.120 8.705 1.260 ;
        RECT 6.575 1.075 6.865 1.120 ;
        RECT 8.415 1.075 8.705 1.120 ;
        RECT 1.470 0.920 1.760 0.965 ;
        RECT 6.990 0.920 7.280 0.965 ;
        RECT 7.910 0.920 8.200 0.965 ;
        RECT 1.470 0.780 8.200 0.920 ;
        RECT 1.470 0.735 1.760 0.780 ;
        RECT 6.990 0.735 7.280 0.780 ;
        RECT 7.910 0.735 8.200 0.780 ;
  END
END sky130_fd_sc_hd__mux4_1

#--------EOF---------

MACRO sky130_fd_sc_hd__mux4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 6.635 1.075 6.945 1.325 ;
        RECT 6.535 0.995 6.945 1.075 ;
        RECT 6.535 0.375 6.845 0.995 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 4.745 0.715 5.115 1.395 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.835 0.765 1.235 1.095 ;
        RECT 1.020 0.395 1.235 0.765 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.410 1.015 2.615 1.320 ;
        RECT 2.240 0.715 2.615 1.015 ;
    END
  END A3
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393000 ;
    PORT
      LAYER met1 ;
        RECT 0.085 1.600 0.375 1.645 ;
        RECT 1.005 1.600 1.295 1.645 ;
        RECT 6.065 1.600 6.355 1.645 ;
        RECT 0.085 1.460 6.355 1.600 ;
        RECT 0.085 1.415 0.375 1.460 ;
        RECT 1.005 1.415 1.295 1.460 ;
        RECT 6.065 1.415 6.355 1.460 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.303000 ;
    PORT
      LAYER li1 ;
        RECT 2.785 0.715 3.075 1.320 ;
    END
  END S1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.825 0.785 8.275 1.015 ;
        RECT 0.005 0.105 8.275 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 7.355 1.835 7.765 2.455 ;
        RECT 7.455 1.495 7.765 1.835 ;
        RECT 7.595 0.725 7.765 1.495 ;
        RECT 7.435 0.265 7.765 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.175 2.085 0.345 2.375 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.410 2.125 2.240 2.295 ;
        RECT 0.175 1.955 0.665 2.085 ;
        RECT 0.175 1.915 1.900 1.955 ;
        RECT 0.495 1.785 1.900 1.915 ;
        RECT 0.145 0.975 0.325 1.745 ;
        RECT 0.495 0.805 0.665 1.785 ;
        RECT 1.005 1.445 1.390 1.615 ;
        RECT 1.220 1.285 1.390 1.445 ;
        RECT 1.560 1.575 1.900 1.785 ;
        RECT 1.560 1.035 1.730 1.575 ;
        RECT 2.070 1.405 2.240 2.125 ;
        RECT 2.595 2.055 2.825 2.635 ;
        RECT 3.305 2.125 3.820 2.295 ;
        RECT 2.970 1.785 3.315 1.955 ;
        RECT 3.565 1.810 3.820 2.125 ;
        RECT 3.145 1.660 3.315 1.785 ;
        RECT 3.145 1.490 3.415 1.660 ;
        RECT 0.170 0.635 0.665 0.805 ;
        RECT 1.405 0.705 1.730 1.035 ;
        RECT 1.900 1.235 2.240 1.405 ;
        RECT 3.245 1.390 3.415 1.490 ;
        RECT 0.170 0.345 0.345 0.635 ;
        RECT 1.900 0.535 2.070 1.235 ;
        RECT 3.245 1.060 3.480 1.390 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.470 0.365 2.070 0.535 ;
        RECT 2.450 0.085 2.780 0.545 ;
        RECT 3.245 0.465 3.415 1.060 ;
        RECT 3.650 0.675 3.820 1.810 ;
        RECT 2.985 0.295 3.415 0.465 ;
        RECT 3.585 0.345 3.820 0.675 ;
        RECT 3.990 2.125 4.515 2.295 ;
        RECT 3.990 0.345 4.180 2.125 ;
        RECT 4.755 2.005 5.100 2.635 ;
        RECT 5.325 2.155 6.275 2.325 ;
        RECT 4.395 1.735 4.585 1.895 ;
        RECT 5.325 1.735 5.495 2.155 ;
        RECT 6.525 2.125 6.845 2.295 ;
        RECT 4.395 1.565 5.495 1.735 ;
        RECT 4.395 0.585 4.565 1.565 ;
        RECT 4.395 0.255 4.600 0.585 ;
        RECT 4.795 0.085 5.125 0.545 ;
        RECT 5.325 0.465 5.495 1.565 ;
        RECT 5.665 1.035 5.955 1.985 ;
        RECT 6.675 1.665 6.845 2.125 ;
        RECT 7.015 1.835 7.185 2.635 ;
        RECT 6.125 1.245 6.465 1.645 ;
        RECT 6.675 1.495 7.285 1.665 ;
        RECT 7.935 1.495 8.185 2.635 ;
        RECT 7.115 1.325 7.285 1.495 ;
        RECT 5.665 0.705 6.285 1.035 ;
        RECT 7.115 0.995 7.425 1.325 ;
        RECT 5.325 0.295 6.220 0.465 ;
        RECT 7.015 0.085 7.265 0.815 ;
        RECT 7.935 0.085 8.190 0.885 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 1.985 2.125 2.155 2.295 ;
        RECT 1.525 1.785 1.695 1.955 ;
        RECT 0.145 1.445 0.315 1.615 ;
        RECT 1.065 1.445 1.235 1.615 ;
        RECT 3.365 2.125 3.535 2.295 ;
        RECT 4.285 2.125 4.455 2.295 ;
        RECT 6.585 2.125 6.755 2.295 ;
        RECT 5.665 1.785 5.835 1.955 ;
        RECT 6.125 1.445 6.295 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
      LAYER met1 ;
        RECT 1.925 2.280 2.215 2.325 ;
        RECT 3.305 2.280 3.595 2.325 ;
        RECT 1.925 2.140 3.595 2.280 ;
        RECT 1.925 2.095 2.215 2.140 ;
        RECT 3.305 2.095 3.595 2.140 ;
        RECT 4.225 2.280 4.515 2.325 ;
        RECT 6.525 2.280 6.815 2.325 ;
        RECT 4.225 2.140 6.815 2.280 ;
        RECT 4.225 2.095 4.515 2.140 ;
        RECT 6.525 2.095 6.815 2.140 ;
        RECT 1.465 1.940 1.755 1.985 ;
        RECT 5.605 1.940 5.895 1.985 ;
        RECT 1.465 1.800 5.895 1.940 ;
        RECT 1.465 1.755 1.755 1.800 ;
        RECT 5.605 1.755 5.895 1.800 ;
  END
END sky130_fd_sc_hd__mux4_2

#--------EOF---------

MACRO sky130_fd_sc_hd__mux4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__mux4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 6.640 1.075 6.950 1.325 ;
        RECT 6.540 0.995 6.950 1.075 ;
        RECT 6.540 0.375 6.850 0.995 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 4.750 0.715 5.120 1.395 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.840 0.765 1.240 1.095 ;
        RECT 1.025 0.395 1.240 0.765 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.415 1.015 2.620 1.320 ;
        RECT 2.245 0.715 2.620 1.015 ;
    END
  END A3
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393000 ;
    PORT
      LAYER met1 ;
        RECT 0.085 1.600 0.380 1.645 ;
        RECT 1.010 1.600 1.300 1.645 ;
        RECT 6.070 1.600 6.360 1.645 ;
        RECT 0.085 1.460 6.360 1.600 ;
        RECT 0.085 1.415 0.380 1.460 ;
        RECT 1.010 1.415 1.300 1.460 ;
        RECT 6.070 1.415 6.360 1.460 ;
    END
  END S0
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.303000 ;
    PORT
      LAYER li1 ;
        RECT 2.790 0.715 3.080 1.320 ;
    END
  END S1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 6.830 0.785 9.195 1.015 ;
        RECT 0.005 0.105 9.195 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.390 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 7.360 1.835 7.770 2.455 ;
        RECT 7.460 1.495 7.770 1.835 ;
        RECT 7.600 1.305 7.770 1.495 ;
        RECT 8.360 1.305 8.685 2.455 ;
        RECT 7.600 1.065 8.685 1.305 ;
        RECT 7.600 0.725 7.770 1.065 ;
        RECT 7.440 0.265 7.770 0.725 ;
        RECT 8.360 0.265 8.685 1.065 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.135 2.085 0.345 2.375 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.415 2.125 2.245 2.295 ;
        RECT 0.135 1.955 0.670 2.085 ;
        RECT 0.135 1.915 1.905 1.955 ;
        RECT 0.500 1.785 1.905 1.915 ;
        RECT 0.150 0.975 0.330 1.745 ;
        RECT 0.500 0.805 0.670 1.785 ;
        RECT 1.010 1.445 1.395 1.615 ;
        RECT 1.225 1.285 1.395 1.445 ;
        RECT 1.565 1.575 1.905 1.785 ;
        RECT 1.565 1.035 1.735 1.575 ;
        RECT 2.075 1.405 2.245 2.125 ;
        RECT 2.600 2.055 2.830 2.635 ;
        RECT 3.310 2.125 3.825 2.295 ;
        RECT 2.975 1.785 3.320 1.955 ;
        RECT 3.575 1.810 3.825 2.125 ;
        RECT 3.150 1.660 3.320 1.785 ;
        RECT 3.150 1.490 3.420 1.660 ;
        RECT 0.135 0.635 0.670 0.805 ;
        RECT 1.410 0.705 1.735 1.035 ;
        RECT 1.905 1.235 2.245 1.405 ;
        RECT 3.250 1.390 3.420 1.490 ;
        RECT 0.135 0.345 0.345 0.635 ;
        RECT 1.905 0.535 2.075 1.235 ;
        RECT 3.250 1.060 3.485 1.390 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.475 0.365 2.075 0.535 ;
        RECT 2.455 0.085 2.785 0.545 ;
        RECT 3.250 0.465 3.420 1.060 ;
        RECT 3.655 0.675 3.825 1.810 ;
        RECT 2.990 0.295 3.420 0.465 ;
        RECT 3.590 0.345 3.825 0.675 ;
        RECT 3.995 2.125 4.520 2.295 ;
        RECT 3.995 0.345 4.185 2.125 ;
        RECT 4.760 2.005 5.105 2.635 ;
        RECT 5.330 2.155 6.280 2.325 ;
        RECT 4.400 1.735 4.590 1.895 ;
        RECT 5.330 1.735 5.500 2.155 ;
        RECT 6.530 2.125 6.850 2.295 ;
        RECT 4.400 1.565 5.500 1.735 ;
        RECT 4.400 0.585 4.570 1.565 ;
        RECT 4.400 0.255 4.605 0.585 ;
        RECT 4.800 0.085 5.130 0.545 ;
        RECT 5.330 0.465 5.500 1.565 ;
        RECT 5.670 1.035 5.960 1.985 ;
        RECT 6.680 1.665 6.850 2.125 ;
        RECT 7.020 1.835 7.190 2.635 ;
        RECT 6.130 1.245 6.470 1.645 ;
        RECT 6.680 1.495 7.290 1.665 ;
        RECT 7.940 1.495 8.190 2.635 ;
        RECT 8.855 1.495 9.105 2.635 ;
        RECT 7.120 1.325 7.290 1.495 ;
        RECT 5.670 0.705 6.290 1.035 ;
        RECT 7.120 0.995 7.430 1.325 ;
        RECT 5.330 0.295 6.225 0.465 ;
        RECT 7.020 0.085 7.270 0.815 ;
        RECT 7.940 0.085 8.190 0.885 ;
        RECT 8.855 0.085 9.105 0.885 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 1.990 2.125 2.160 2.295 ;
        RECT 1.530 1.785 1.700 1.955 ;
        RECT 0.150 1.445 0.320 1.615 ;
        RECT 1.070 1.445 1.240 1.615 ;
        RECT 3.370 2.125 3.540 2.295 ;
        RECT 4.290 2.125 4.460 2.295 ;
        RECT 6.590 2.125 6.760 2.295 ;
        RECT 5.670 1.785 5.840 1.955 ;
        RECT 6.130 1.445 6.300 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
      LAYER met1 ;
        RECT 1.930 2.280 2.220 2.325 ;
        RECT 3.310 2.280 3.600 2.325 ;
        RECT 1.930 2.140 3.600 2.280 ;
        RECT 1.930 2.095 2.220 2.140 ;
        RECT 3.310 2.095 3.600 2.140 ;
        RECT 4.230 2.280 4.520 2.325 ;
        RECT 6.530 2.280 6.820 2.325 ;
        RECT 4.230 2.140 6.820 2.280 ;
        RECT 4.230 2.095 4.520 2.140 ;
        RECT 6.530 2.095 6.820 2.140 ;
        RECT 1.470 1.940 1.760 1.985 ;
        RECT 5.610 1.940 5.900 1.985 ;
        RECT 1.470 1.800 5.900 1.940 ;
        RECT 1.470 1.755 1.760 1.800 ;
        RECT 5.610 1.755 5.900 1.800 ;
  END
END sky130_fd_sc_hd__mux4_4

#--------EOF---------

MACRO sky130_fd_sc_hd__nand2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.940 1.075 1.275 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.055 0.430 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.105 1.375 1.015 ;
        RECT 0.140 -0.085 0.310 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.485 0.865 2.465 ;
        RECT 0.600 0.885 0.770 1.485 ;
        RECT 0.600 0.255 1.295 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.085 1.495 0.365 2.635 ;
        RECT 1.035 1.495 1.295 2.635 ;
        RECT 0.085 0.085 0.395 0.885 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
END sky130_fd_sc_hd__nand2_1

#--------EOF---------

MACRO sky130_fd_sc_hd__nand2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.075 1.765 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.845 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.195 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.715500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 0.515 1.495 2.215 1.665 ;
        RECT 1.935 0.905 2.215 1.495 ;
        RECT 1.355 0.655 2.215 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.110 2.635 ;
        RECT 0.085 0.715 1.185 0.885 ;
        RECT 0.085 0.255 0.425 0.715 ;
        RECT 0.595 0.085 0.765 0.545 ;
        RECT 0.935 0.465 1.185 0.715 ;
        RECT 1.775 0.465 2.105 0.485 ;
        RECT 0.935 0.255 2.105 0.465 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__nand2_2

#--------EOF---------

MACRO sky130_fd_sc_hd__nand2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 2.615 1.075 4.055 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 1.730 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.875 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.431000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.195 1.665 2.525 2.465 ;
        RECT 3.035 1.665 3.365 2.465 ;
        RECT 0.515 1.495 3.365 1.665 ;
        RECT 1.910 1.075 2.445 1.495 ;
        RECT 2.195 0.805 2.445 1.075 ;
        RECT 2.195 0.635 3.365 0.805 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.025 2.635 ;
        RECT 2.695 1.835 2.865 2.635 ;
        RECT 3.535 1.835 3.785 2.635 ;
        RECT 0.090 0.715 2.025 0.905 ;
        RECT 0.090 0.255 0.425 0.715 ;
        RECT 0.595 0.085 0.765 0.545 ;
        RECT 0.935 0.255 1.265 0.715 ;
        RECT 1.435 0.085 1.605 0.545 ;
        RECT 1.775 0.465 2.025 0.715 ;
        RECT 3.535 0.465 3.785 0.885 ;
        RECT 1.775 0.255 3.785 0.465 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__nand2_4

#--------EOF---------

MACRO sky130_fd_sc_hd__nand2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 4.290 1.075 6.305 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 0.510 1.075 3.365 1.295 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.355 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.862000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.195 1.665 2.525 2.465 ;
        RECT 3.035 1.665 3.365 2.465 ;
        RECT 3.875 1.665 4.205 2.465 ;
        RECT 4.715 1.665 5.045 2.465 ;
        RECT 5.555 1.665 5.885 2.465 ;
        RECT 6.395 1.665 6.725 2.465 ;
        RECT 0.515 1.465 6.725 1.665 ;
        RECT 3.640 1.075 4.120 1.465 ;
        RECT 3.875 0.905 4.120 1.075 ;
        RECT 6.475 0.905 6.725 1.465 ;
        RECT 3.875 0.655 6.725 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.025 2.635 ;
        RECT 2.695 1.835 2.865 2.635 ;
        RECT 3.535 1.835 3.705 2.635 ;
        RECT 4.375 1.835 4.545 2.635 ;
        RECT 5.215 1.835 5.385 2.635 ;
        RECT 6.055 1.835 6.225 2.635 ;
        RECT 6.915 1.495 7.270 2.635 ;
        RECT 0.090 0.735 3.705 0.905 ;
        RECT 0.090 0.255 0.425 0.735 ;
        RECT 0.595 0.085 0.765 0.565 ;
        RECT 0.935 0.255 1.265 0.735 ;
        RECT 1.435 0.085 1.605 0.565 ;
        RECT 1.775 0.255 2.105 0.735 ;
        RECT 2.275 0.085 2.445 0.565 ;
        RECT 2.615 0.255 2.945 0.735 ;
        RECT 3.115 0.085 3.285 0.565 ;
        RECT 3.455 0.485 3.705 0.735 ;
        RECT 6.895 0.485 7.270 0.905 ;
        RECT 3.455 0.255 7.270 0.485 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
END sky130_fd_sc_hd__nand2_8

#--------EOF---------

MACRO sky130_fd_sc_hd__nand2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.440 1.315 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.610 1.075 1.085 1.315 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 1.840 1.015 ;
        RECT 0.150 0.105 1.840 0.335 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 1.000 2.005 1.330 2.465 ;
        RECT 1.000 1.835 2.170 2.005 ;
        RECT 1.800 0.545 2.170 1.835 ;
        RECT 1.420 0.255 2.170 0.545 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.580 1.835 0.830 2.635 ;
        RECT 1.500 2.175 1.715 2.635 ;
        RECT 0.090 1.665 0.370 1.825 ;
        RECT 0.090 1.495 1.425 1.665 ;
        RECT 1.255 1.325 1.425 1.495 ;
        RECT 1.255 1.075 1.630 1.325 ;
        RECT 1.255 0.905 1.425 1.075 ;
        RECT 0.090 0.735 1.425 0.905 ;
        RECT 0.090 0.525 0.360 0.735 ;
        RECT 0.580 0.085 0.910 0.545 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__nand2b_1

#--------EOF---------

MACRO sky130_fd_sc_hd__nand2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.455 0.995 0.800 1.325 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.990 1.275 2.180 1.655 ;
        RECT 1.990 1.075 3.135 1.275 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 3.205 1.015 ;
        RECT 0.150 0.105 3.205 0.335 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.775500 ;
    PORT
      LAYER li1 ;
        RECT 1.035 2.005 1.365 2.465 ;
        RECT 2.280 2.005 2.635 2.465 ;
        RECT 1.035 1.835 2.635 2.005 ;
        RECT 1.530 0.905 1.810 1.835 ;
        RECT 2.360 1.495 2.635 1.835 ;
        RECT 1.530 0.805 1.855 0.905 ;
        RECT 1.525 0.635 1.855 0.805 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.110 1.665 0.410 1.860 ;
        RECT 0.580 1.835 0.835 2.635 ;
        RECT 1.535 2.175 2.110 2.635 ;
        RECT 0.110 1.495 1.360 1.665 ;
        RECT 2.805 1.495 3.135 2.635 ;
        RECT 0.110 0.840 0.280 1.495 ;
        RECT 1.030 1.075 1.360 1.495 ;
        RECT 0.110 0.510 0.345 0.840 ;
        RECT 0.515 0.085 0.845 0.825 ;
        RECT 1.080 0.465 1.355 0.905 ;
        RECT 2.025 0.695 3.135 0.905 ;
        RECT 2.025 0.465 2.275 0.695 ;
        RECT 1.080 0.255 2.275 0.465 ;
        RECT 2.445 0.085 2.615 0.525 ;
        RECT 2.785 0.255 3.135 0.695 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__nand2b_2

#--------EOF---------

MACRO sky130_fd_sc_hd__nand2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand2b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.440 1.275 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.155 1.075 4.940 1.275 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.960 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.431000 ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.665 1.785 2.465 ;
        RECT 2.295 1.665 2.640 2.465 ;
        RECT 3.150 1.665 3.480 2.465 ;
        RECT 3.990 1.665 4.320 2.465 ;
        RECT 1.455 1.445 4.320 1.665 ;
        RECT 2.375 0.905 2.640 1.445 ;
        RECT 1.455 0.635 2.640 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.090 1.665 0.425 2.465 ;
        RECT 0.595 1.835 1.285 2.635 ;
        RECT 1.955 1.835 2.125 2.635 ;
        RECT 2.810 1.835 2.980 2.635 ;
        RECT 3.650 1.835 3.820 2.635 ;
        RECT 0.090 1.445 0.780 1.665 ;
        RECT 0.970 1.445 1.285 1.835 ;
        RECT 4.520 1.495 4.850 2.635 ;
        RECT 0.610 1.275 0.780 1.445 ;
        RECT 0.610 1.075 2.205 1.275 ;
        RECT 0.610 0.905 0.780 1.075 ;
        RECT 0.090 0.715 0.780 0.905 ;
        RECT 0.090 0.255 0.425 0.715 ;
        RECT 0.595 0.085 0.790 0.545 ;
        RECT 1.035 0.465 1.285 0.905 ;
        RECT 2.810 0.715 4.850 0.905 ;
        RECT 2.810 0.465 3.060 0.715 ;
        RECT 1.035 0.255 3.060 0.465 ;
        RECT 3.230 0.085 3.400 0.545 ;
        RECT 3.570 0.255 3.900 0.715 ;
        RECT 4.070 0.085 4.310 0.545 ;
        RECT 4.520 0.255 4.850 0.715 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
END sky130_fd_sc_hd__nand2b_4

#--------EOF---------

MACRO sky130_fd_sc_hd__nand3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.445 0.995 1.755 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.865 0.765 1.240 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 0.745 0.330 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.835 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.699000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.415 1.665 1.745 2.465 ;
        RECT 0.515 1.495 1.745 1.665 ;
        RECT 0.515 0.595 0.695 1.495 ;
        RECT 1.415 0.595 1.745 0.825 ;
        RECT 0.515 0.255 1.745 0.595 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.245 2.635 ;
        RECT 0.090 0.085 0.345 0.575 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__nand3_1

#--------EOF---------

MACRO sky130_fd_sc_hd__nand3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.995 0.330 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.070 1.075 2.160 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.470 1.075 3.595 1.275 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.605 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.985500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.715 1.665 3.045 2.465 ;
        RECT 0.515 1.445 3.045 1.665 ;
        RECT 0.515 0.635 0.845 1.445 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.545 2.635 ;
        RECT 3.215 1.445 3.595 2.635 ;
        RECT 0.090 0.465 0.345 0.785 ;
        RECT 1.355 0.635 3.045 0.905 ;
        RECT 0.090 0.295 2.105 0.465 ;
        RECT 2.295 0.085 2.625 0.465 ;
        RECT 3.215 0.085 3.595 0.885 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__nand3_2

#--------EOF---------

MACRO sky130_fd_sc_hd__nand3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.850 1.075 5.565 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.990 1.075 3.540 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 1.700 1.275 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.085 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.971000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.195 1.665 2.525 2.465 ;
        RECT 3.035 1.665 3.365 2.465 ;
        RECT 4.395 1.665 4.725 2.465 ;
        RECT 5.235 1.665 5.565 2.465 ;
        RECT 0.515 1.445 6.355 1.665 ;
        RECT 6.125 0.905 6.355 1.445 ;
        RECT 4.395 0.655 6.355 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.090 1.445 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.025 2.635 ;
        RECT 2.695 1.835 2.865 2.635 ;
        RECT 3.535 1.835 4.225 2.635 ;
        RECT 4.895 1.835 5.065 2.635 ;
        RECT 5.735 1.835 6.000 2.635 ;
        RECT 0.090 0.735 3.785 0.905 ;
        RECT 0.090 0.255 0.425 0.735 ;
        RECT 0.595 0.085 0.765 0.565 ;
        RECT 0.935 0.255 1.265 0.735 ;
        RECT 1.775 0.655 2.105 0.735 ;
        RECT 2.615 0.655 2.945 0.735 ;
        RECT 3.455 0.655 3.785 0.735 ;
        RECT 1.435 0.085 1.605 0.565 ;
        RECT 2.195 0.255 6.000 0.485 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
END sky130_fd_sc_hd__nand3_4

#--------EOF---------

MACRO sky130_fd_sc_hd__nand3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.325 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.425 0.995 1.755 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.965 0.995 1.235 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.135 0.335 2.525 1.015 ;
        RECT 0.145 0.105 2.525 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.732000 ;
    PORT
      LAYER li1 ;
        RECT 1.130 1.665 1.460 2.465 ;
        RECT 2.085 1.665 2.675 2.465 ;
        RECT 1.130 1.495 2.675 1.665 ;
        RECT 2.385 0.485 2.675 1.495 ;
        RECT 2.085 0.255 2.675 0.485 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.085 1.595 0.510 1.925 ;
        RECT 0.085 0.825 0.255 1.595 ;
        RECT 0.710 1.495 0.960 2.635 ;
        RECT 1.630 1.835 1.915 2.635 ;
        RECT 2.045 0.825 2.215 1.325 ;
        RECT 0.085 0.655 2.215 0.825 ;
        RECT 0.085 0.445 0.510 0.655 ;
        RECT 0.710 0.085 1.040 0.485 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__nand3b_1

#--------EOF---------

MACRO sky130_fd_sc_hd__nand3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.430 1.075 0.780 1.275 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.950 1.075 3.140 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.060 1.075 1.740 1.275 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.490 0.785 4.100 1.015 ;
        RECT 0.005 0.105 4.100 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.985500 ;
    PORT
      LAYER li1 ;
        RECT 1.060 2.005 1.390 2.465 ;
        RECT 1.900 2.005 2.230 2.465 ;
        RECT 1.060 1.955 2.230 2.005 ;
        RECT 3.260 2.005 3.510 2.465 ;
        RECT 3.260 1.955 4.050 2.005 ;
        RECT 1.060 1.785 4.050 1.955 ;
        RECT 3.850 0.905 4.050 1.785 ;
        RECT 3.260 0.635 4.050 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.090 2.065 0.410 2.465 ;
        RECT 0.090 1.615 0.260 2.065 ;
        RECT 0.580 1.835 0.890 2.635 ;
        RECT 1.560 2.175 1.730 2.635 ;
        RECT 2.400 2.175 2.650 2.635 ;
        RECT 2.840 2.175 3.090 2.635 ;
        RECT 3.760 2.175 4.050 2.635 ;
        RECT 0.090 1.445 3.650 1.615 ;
        RECT 0.090 0.655 0.260 1.445 ;
        RECT 3.320 1.075 3.650 1.445 ;
        RECT 0.090 0.255 0.410 0.655 ;
        RECT 0.580 0.085 0.890 0.905 ;
        RECT 1.060 0.715 2.750 0.905 ;
        RECT 1.060 0.255 1.390 0.715 ;
        RECT 2.000 0.635 2.750 0.715 ;
        RECT 1.560 0.085 1.810 0.545 ;
        RECT 2.920 0.465 3.090 0.905 ;
        RECT 2.000 0.255 4.050 0.465 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__nand3b_2

#--------EOF---------

MACRO sky130_fd_sc_hd__nand3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand3b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.430 1.075 0.780 1.275 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.270 1.075 4.480 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 4.790 1.075 6.500 1.275 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.115 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.971000 ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.665 1.785 2.465 ;
        RECT 2.295 2.005 2.625 2.465 ;
        RECT 3.135 2.005 3.465 2.465 ;
        RECT 2.295 1.665 3.465 2.005 ;
        RECT 3.975 1.665 4.305 2.465 ;
        RECT 5.335 1.665 5.665 2.465 ;
        RECT 6.175 1.665 6.505 2.465 ;
        RECT 1.455 1.445 6.505 1.665 ;
        RECT 2.795 1.075 3.100 1.445 ;
        RECT 2.795 0.905 2.965 1.075 ;
        RECT 1.455 0.635 2.965 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.085 1.445 0.425 2.465 ;
        RECT 0.595 1.445 1.285 2.635 ;
        RECT 1.955 1.835 2.125 2.635 ;
        RECT 2.795 2.175 2.965 2.635 ;
        RECT 3.635 1.835 3.805 2.635 ;
        RECT 4.475 1.835 5.165 2.635 ;
        RECT 5.835 1.835 6.005 2.635 ;
        RECT 6.675 1.445 7.005 2.635 ;
        RECT 0.085 0.905 0.260 1.445 ;
        RECT 1.005 1.075 2.625 1.275 ;
        RECT 1.005 0.905 1.285 1.075 ;
        RECT 0.085 0.715 1.285 0.905 ;
        RECT 3.135 0.715 6.505 0.905 ;
        RECT 0.085 0.255 0.425 0.715 ;
        RECT 3.135 0.635 4.725 0.715 ;
        RECT 0.595 0.085 0.845 0.545 ;
        RECT 1.035 0.255 4.725 0.465 ;
        RECT 4.915 0.085 5.165 0.545 ;
        RECT 5.335 0.255 5.665 0.715 ;
        RECT 5.835 0.085 6.005 0.545 ;
        RECT 6.175 0.255 6.505 0.715 ;
        RECT 6.675 0.085 7.005 0.905 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
END sky130_fd_sc_hd__nand3b_4

#--------EOF---------

MACRO sky130_fd_sc_hd__nand4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.975 0.995 2.215 1.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.145 0.995 1.455 1.325 ;
        RECT 1.145 0.825 1.350 0.995 ;
        RECT 1.000 0.300 1.350 0.825 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.995 0.975 1.325 ;
        RECT 0.595 0.300 0.810 0.995 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 0.995 0.395 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.295 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.385 1.665 1.715 2.465 ;
        RECT 0.515 1.495 1.795 1.665 ;
        RECT 1.625 0.825 1.795 1.495 ;
        RECT 1.520 0.255 2.215 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.915 1.835 2.195 2.635 ;
        RECT 0.090 0.085 0.425 0.825 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__nand4_1

#--------EOF---------

MACRO sky130_fd_sc_hd__nand4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.165 1.075 4.495 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.235 1.075 3.080 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.070 1.075 1.700 1.275 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.845 1.275 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.535 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.255500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.355 1.665 2.685 2.465 ;
        RECT 3.595 1.665 3.925 2.465 ;
        RECT 0.515 1.445 3.925 1.665 ;
        RECT 3.370 1.055 3.925 1.445 ;
        RECT 3.595 0.635 3.925 1.055 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.185 2.635 ;
        RECT 2.995 1.835 3.325 2.635 ;
        RECT 4.095 1.445 4.425 2.635 ;
        RECT 0.090 0.735 1.185 0.905 ;
        RECT 0.090 0.255 0.425 0.735 ;
        RECT 0.595 0.085 0.765 0.545 ;
        RECT 0.935 0.465 1.185 0.735 ;
        RECT 1.355 0.635 3.085 0.905 ;
        RECT 3.255 0.465 3.425 0.885 ;
        RECT 4.095 0.465 4.425 0.905 ;
        RECT 0.935 0.255 2.125 0.465 ;
        RECT 2.315 0.255 4.425 0.465 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__nand4_2

#--------EOF---------

MACRO sky130_fd_sc_hd__nand4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.465 1.075 7.710 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.850 1.075 5.565 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.990 1.075 3.540 1.275 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 1.700 1.275 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.815 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.511000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 2.195 1.665 2.525 2.465 ;
        RECT 3.035 1.665 3.365 2.465 ;
        RECT 4.395 1.665 4.725 2.465 ;
        RECT 5.235 1.665 5.565 2.465 ;
        RECT 6.135 1.665 6.465 2.465 ;
        RECT 6.975 1.665 7.305 2.465 ;
        RECT 0.515 1.445 7.305 1.665 ;
        RECT 6.110 0.905 6.290 1.445 ;
        RECT 6.110 0.655 7.305 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.090 1.445 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.025 2.635 ;
        RECT 2.695 1.835 2.865 2.635 ;
        RECT 3.535 1.835 4.225 2.635 ;
        RECT 4.895 1.835 5.065 2.635 ;
        RECT 5.770 1.835 5.940 2.635 ;
        RECT 6.635 1.835 6.805 2.635 ;
        RECT 7.475 1.445 7.735 2.635 ;
        RECT 0.090 0.655 2.025 0.905 ;
        RECT 2.195 0.655 5.565 0.905 ;
        RECT 0.090 0.255 0.345 0.655 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.015 0.255 1.185 0.655 ;
        RECT 1.855 0.485 2.025 0.655 ;
        RECT 5.770 0.485 5.940 0.905 ;
        RECT 7.475 0.485 7.730 0.905 ;
        RECT 1.355 0.085 1.685 0.485 ;
        RECT 1.855 0.255 3.785 0.485 ;
        RECT 3.975 0.255 7.730 0.485 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
  END
END sky130_fd_sc_hd__nand4_4

#--------EOF---------

MACRO sky130_fd_sc_hd__nand4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.325 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.925 0.765 2.185 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.505 0.765 1.755 1.325 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.965 0.995 1.235 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.075 0.335 3.135 1.015 ;
        RECT 0.145 0.105 3.135 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.887500 ;
    PORT
      LAYER li1 ;
        RECT 1.130 1.665 1.460 2.465 ;
        RECT 2.085 1.665 2.415 2.465 ;
        RECT 1.130 1.495 3.135 1.665 ;
        RECT 2.925 0.825 3.135 1.495 ;
        RECT 2.695 0.255 3.135 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.595 0.510 1.925 ;
        RECT 0.085 0.825 0.255 1.595 ;
        RECT 0.710 1.495 0.960 2.635 ;
        RECT 1.630 1.835 1.915 2.635 ;
        RECT 2.705 1.835 2.920 2.635 ;
        RECT 2.355 0.995 2.755 1.325 ;
        RECT 0.085 0.655 1.335 0.825 ;
        RECT 0.085 0.445 0.475 0.655 ;
        RECT 1.155 0.595 1.335 0.655 ;
        RECT 2.355 0.595 2.525 0.995 ;
        RECT 0.655 0.085 0.985 0.485 ;
        RECT 1.155 0.425 2.525 0.595 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__nand4b_1

#--------EOF---------

MACRO sky130_fd_sc_hd__nand4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.995 0.330 1.615 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.010 1.075 3.100 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.360 1.075 4.450 1.275 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.620 1.075 5.430 1.275 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.945 0.785 5.425 1.015 ;
        RECT 0.005 0.105 5.425 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.255500 ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.665 1.785 2.465 ;
        RECT 2.295 1.665 2.625 2.465 ;
        RECT 3.605 1.665 3.935 2.465 ;
        RECT 4.535 1.665 4.865 2.465 ;
        RECT 1.455 1.445 4.865 1.665 ;
        RECT 1.550 0.825 1.785 1.445 ;
        RECT 1.455 0.635 1.785 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.090 2.085 0.345 2.465 ;
        RECT 0.515 2.255 1.285 2.635 ;
        RECT 0.090 1.915 0.670 2.085 ;
        RECT 0.500 1.245 0.670 1.915 ;
        RECT 1.035 1.445 1.285 2.255 ;
        RECT 1.955 1.835 2.125 2.635 ;
        RECT 2.795 1.835 3.435 2.635 ;
        RECT 4.105 1.835 4.365 2.635 ;
        RECT 5.035 1.495 5.430 2.635 ;
        RECT 0.500 1.075 1.380 1.245 ;
        RECT 0.500 0.805 0.670 1.075 ;
        RECT 0.090 0.635 0.670 0.805 ;
        RECT 0.090 0.255 0.345 0.635 ;
        RECT 1.035 0.465 1.285 0.905 ;
        RECT 1.955 0.635 3.045 0.905 ;
        RECT 3.235 0.715 5.340 0.905 ;
        RECT 3.235 0.635 4.455 0.715 ;
        RECT 1.955 0.465 2.125 0.635 ;
        RECT 4.155 0.615 4.455 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.035 0.255 2.125 0.465 ;
        RECT 2.295 0.255 3.985 0.465 ;
        RECT 4.155 0.255 4.415 0.615 ;
        RECT 4.665 0.085 4.835 0.545 ;
        RECT 5.005 0.255 5.340 0.715 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__nand4b_2

#--------EOF---------

MACRO sky130_fd_sc_hd__nand4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.440 1.275 ;
    END
  END A_N
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 2.930 1.075 4.590 1.275 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 4.790 1.075 6.510 1.275 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 7.015 1.075 8.655 1.275 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.695 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.511000 ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.665 1.785 2.465 ;
        RECT 2.295 1.665 2.625 2.465 ;
        RECT 3.135 1.665 3.465 2.465 ;
        RECT 3.975 1.665 4.305 2.465 ;
        RECT 5.335 1.665 5.665 2.465 ;
        RECT 6.175 1.665 6.505 2.465 ;
        RECT 7.015 1.665 7.345 2.465 ;
        RECT 7.855 1.665 8.185 2.465 ;
        RECT 1.455 1.445 8.185 1.665 ;
        RECT 2.375 0.905 2.640 1.445 ;
        RECT 1.455 0.635 2.640 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.740 2.805 ;
        RECT 0.090 1.665 0.425 2.465 ;
        RECT 0.595 1.835 1.285 2.635 ;
        RECT 1.955 1.835 2.125 2.635 ;
        RECT 2.795 1.835 2.965 2.635 ;
        RECT 3.635 1.835 3.805 2.635 ;
        RECT 4.475 1.835 5.165 2.635 ;
        RECT 5.835 1.835 6.005 2.635 ;
        RECT 6.675 1.835 6.845 2.635 ;
        RECT 7.515 1.835 7.685 2.635 ;
        RECT 0.090 1.495 0.805 1.665 ;
        RECT 0.995 1.495 1.285 1.835 ;
        RECT 0.610 1.275 0.805 1.495 ;
        RECT 8.355 1.445 8.610 2.635 ;
        RECT 0.610 1.075 2.205 1.275 ;
        RECT 0.610 0.905 0.805 1.075 ;
        RECT 0.090 0.735 0.805 0.905 ;
        RECT 0.090 0.255 0.425 0.735 ;
        RECT 0.595 0.085 0.845 0.545 ;
        RECT 1.035 0.465 1.285 0.905 ;
        RECT 3.135 0.635 6.505 0.905 ;
        RECT 6.675 0.735 8.610 0.905 ;
        RECT 6.675 0.465 6.925 0.735 ;
        RECT 1.035 0.255 4.725 0.465 ;
        RECT 4.915 0.255 6.925 0.465 ;
        RECT 7.095 0.085 7.265 0.545 ;
        RECT 7.435 0.255 7.765 0.735 ;
        RECT 7.935 0.085 8.105 0.545 ;
        RECT 8.275 0.255 8.610 0.735 ;
        RECT 0.000 -0.085 8.740 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
  END
END sky130_fd_sc_hd__nand4b_4

#--------EOF---------

MACRO sky130_fd_sc_hd__nand4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4bb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 3.390 0.725 3.640 1.615 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.430 1.075 0.780 1.655 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.500 0.735 1.720 1.325 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.970 1.075 1.320 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 3.020 1.015 ;
        RECT 0.005 0.335 4.135 0.785 ;
        RECT 0.145 0.105 4.135 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.909000 ;
    PORT
      LAYER li1 ;
        RECT 1.120 1.665 1.450 2.465 ;
        RECT 2.140 1.665 2.470 2.465 ;
        RECT 1.120 1.495 2.670 1.665 ;
        RECT 2.420 0.825 2.670 1.495 ;
        RECT 2.420 0.255 2.930 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 2.065 0.425 2.465 ;
        RECT 0.085 0.905 0.260 2.065 ;
        RECT 0.595 1.835 0.925 2.635 ;
        RECT 1.640 1.835 1.970 2.635 ;
        RECT 2.680 2.175 3.450 2.635 ;
        RECT 3.635 2.005 4.055 2.465 ;
        RECT 2.840 1.835 4.055 2.005 ;
        RECT 0.085 0.715 1.270 0.905 ;
        RECT 0.085 0.485 0.425 0.715 ;
        RECT 1.080 0.555 1.270 0.715 ;
        RECT 1.970 0.555 2.250 1.325 ;
        RECT 2.840 0.995 3.090 1.835 ;
        RECT 0.595 0.085 0.900 0.545 ;
        RECT 1.080 0.365 2.250 0.555 ;
        RECT 3.810 0.545 4.055 1.835 ;
        RECT 3.100 0.085 3.450 0.545 ;
        RECT 3.620 0.255 4.055 0.545 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__nand4bb_1

#--------EOF---------

MACRO sky130_fd_sc_hd__nand4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4bb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.610 1.340 0.890 1.615 ;
        RECT 0.560 1.170 0.890 1.340 ;
        RECT 0.610 1.070 0.890 1.170 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.070 0.330 1.615 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.720 1.075 4.615 1.275 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.945 1.075 5.875 1.275 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.575 0.785 5.965 1.015 ;
        RECT 0.005 0.105 5.965 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.255500 ;
    PORT
      LAYER li1 ;
        RECT 2.085 1.665 2.335 2.465 ;
        RECT 2.925 1.665 3.255 2.465 ;
        RECT 4.285 1.665 4.615 2.465 ;
        RECT 5.125 1.665 5.455 2.465 ;
        RECT 2.085 1.445 5.455 1.665 ;
        RECT 2.085 0.655 2.415 1.445 ;
        RECT 3.245 1.075 3.550 1.445 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.085 1.980 0.370 2.440 ;
        RECT 0.540 2.195 0.765 2.635 ;
        RECT 0.935 2.150 1.575 2.465 ;
        RECT 0.085 1.785 1.230 1.980 ;
        RECT 1.060 0.900 1.230 1.785 ;
        RECT 0.085 0.730 1.230 0.900 ;
        RECT 1.400 1.410 1.575 2.150 ;
        RECT 1.745 1.495 1.915 2.635 ;
        RECT 2.505 1.835 2.755 2.635 ;
        RECT 3.425 1.835 4.115 2.635 ;
        RECT 4.785 1.835 4.955 2.635 ;
        RECT 5.625 1.445 5.895 2.635 ;
        RECT 0.085 0.255 0.345 0.730 ;
        RECT 1.400 0.715 1.580 1.410 ;
        RECT 2.745 1.075 3.075 1.275 ;
        RECT 1.400 0.560 1.575 0.715 ;
        RECT 2.925 0.655 4.615 0.905 ;
        RECT 4.785 0.735 5.895 0.905 ;
        RECT 0.515 0.085 0.765 0.545 ;
        RECT 0.935 0.255 1.575 0.560 ;
        RECT 1.745 0.485 1.915 0.585 ;
        RECT 4.785 0.485 5.035 0.735 ;
        RECT 1.745 0.255 3.675 0.485 ;
        RECT 3.865 0.255 5.035 0.485 ;
        RECT 5.205 0.085 5.375 0.565 ;
        RECT 5.545 0.255 5.895 0.735 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 1.060 1.105 1.230 1.275 ;
        RECT 2.905 1.105 3.075 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
      LAYER met1 ;
        RECT 1.000 1.075 3.135 1.305 ;
  END
END sky130_fd_sc_hd__nand4bb_2

#--------EOF---------

MACRO sky130_fd_sc_hd__nand4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nand4bb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.100 0.995 0.330 1.615 ;
    END
  END A_N
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.590 0.995 0.975 1.615 ;
    END
  END B_N
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.120 1.075 7.910 1.275 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 8.420 1.075 10.015 1.275 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 10.115 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.511000 ;
    PORT
      LAYER li1 ;
        RECT 2.540 1.665 2.790 2.465 ;
        RECT 3.380 1.665 3.710 2.465 ;
        RECT 4.220 1.665 4.550 2.465 ;
        RECT 5.060 1.665 5.390 2.465 ;
        RECT 6.740 1.665 7.070 2.465 ;
        RECT 7.580 1.665 7.910 2.465 ;
        RECT 8.420 1.665 8.750 2.465 ;
        RECT 9.260 1.665 9.590 2.465 ;
        RECT 2.540 1.445 9.590 1.665 ;
        RECT 3.700 0.905 3.990 1.445 ;
        RECT 2.540 0.655 3.990 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.085 1.980 0.370 2.440 ;
        RECT 0.540 2.195 0.765 2.635 ;
        RECT 0.935 2.150 1.795 2.465 ;
        RECT 0.085 1.785 1.455 1.980 ;
        RECT 1.145 0.805 1.455 1.785 ;
        RECT 0.085 0.635 1.455 0.805 ;
        RECT 1.625 1.305 1.795 2.150 ;
        RECT 2.200 1.495 2.370 2.635 ;
        RECT 2.960 1.835 3.210 2.635 ;
        RECT 3.880 1.835 4.050 2.635 ;
        RECT 4.720 1.835 4.890 2.635 ;
        RECT 5.610 1.835 6.540 2.635 ;
        RECT 7.240 1.835 7.410 2.635 ;
        RECT 8.080 1.835 8.250 2.635 ;
        RECT 8.920 1.835 9.090 2.635 ;
        RECT 9.760 1.445 10.035 2.635 ;
        RECT 1.625 1.075 2.210 1.305 ;
        RECT 2.540 1.075 3.285 1.245 ;
        RECT 4.160 1.075 5.390 1.275 ;
        RECT 0.085 0.255 0.345 0.635 ;
        RECT 1.625 0.465 1.795 1.075 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.255 1.795 0.465 ;
        RECT 2.200 0.485 2.370 0.905 ;
        RECT 4.220 0.735 6.150 0.905 ;
        RECT 4.220 0.655 5.390 0.735 ;
        RECT 5.980 0.485 6.150 0.735 ;
        RECT 6.320 0.655 10.035 0.905 ;
        RECT 2.200 0.255 5.810 0.485 ;
        RECT 5.980 0.255 7.910 0.485 ;
        RECT 8.420 0.085 8.750 0.485 ;
        RECT 9.260 0.085 9.590 0.485 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 1.980 1.105 2.150 1.275 ;
        RECT 4.280 1.105 4.450 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
      LAYER met1 ;
        RECT 1.920 1.260 2.210 1.305 ;
        RECT 4.220 1.260 4.510 1.305 ;
        RECT 1.920 1.120 4.510 1.260 ;
        RECT 1.920 1.075 2.210 1.120 ;
        RECT 4.220 1.075 4.510 1.120 ;
  END
END sky130_fd_sc_hd__nand4bb_4

#--------EOF---------

MACRO sky130_fd_sc_hd__nor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.380 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.075 1.295 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.435 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.380 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.355 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.570 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.380 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.435500 ;
    PORT
      LAYER li1 ;
        RECT 0.095 1.665 0.425 2.450 ;
        RECT 0.095 1.495 0.775 1.665 ;
        RECT 0.605 0.895 0.775 1.495 ;
        RECT 0.515 0.255 0.845 0.895 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.380 2.805 ;
        RECT 0.955 1.495 1.285 2.635 ;
        RECT 0.105 0.085 0.345 0.895 ;
        RECT 1.015 0.085 1.285 0.895 ;
        RECT 0.000 -0.085 1.380 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
  END
END sky130_fd_sc_hd__nor2_1

#--------EOF---------

MACRO sky130_fd_sc_hd__nor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.810 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.980 1.075 1.750 1.275 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.215 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.621000 ;
    PORT
      LAYER li1 ;
        RECT 1.375 1.665 1.705 2.125 ;
        RECT 1.375 1.445 2.135 1.665 ;
        RECT 1.920 0.905 2.135 1.445 ;
        RECT 0.535 0.735 2.135 0.905 ;
        RECT 0.535 0.725 1.705 0.735 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 1.375 0.255 1.705 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.090 1.665 0.365 2.465 ;
        RECT 0.535 1.835 0.865 2.635 ;
        RECT 1.035 2.295 2.175 2.465 ;
        RECT 1.035 1.665 1.205 2.295 ;
        RECT 1.875 1.835 2.175 2.295 ;
        RECT 0.090 1.455 1.205 1.665 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.165 0.555 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__nor2_2

#--------EOF---------

MACRO sky130_fd_sc_hd__nor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.140 1.075 1.800 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 2.120 1.075 3.485 1.275 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.895 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER li1 ;
        RECT 2.295 1.745 2.465 2.125 ;
        RECT 3.135 1.745 3.305 2.125 ;
        RECT 2.295 1.445 4.055 1.745 ;
        RECT 3.655 0.905 4.055 1.445 ;
        RECT 0.535 0.725 4.055 0.905 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 3.055 0.255 3.385 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.090 1.665 0.365 2.465 ;
        RECT 0.535 1.835 0.865 2.635 ;
        RECT 1.035 1.665 1.205 2.465 ;
        RECT 1.375 1.835 1.625 2.635 ;
        RECT 1.795 2.295 3.890 2.465 ;
        RECT 1.795 1.665 2.125 2.295 ;
        RECT 2.635 1.935 2.965 2.295 ;
        RECT 3.475 1.915 3.890 2.295 ;
        RECT 0.090 1.455 2.125 1.665 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.555 ;
        RECT 2.715 0.085 2.885 0.555 ;
        RECT 3.555 0.085 3.840 0.555 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__nor2_4

#--------EOF---------

MACRO sky130_fd_sc_hd__nor2_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 0.360 1.075 3.530 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 3.800 1.075 6.540 1.275 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.255 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.484000 ;
    PORT
      LAYER li1 ;
        RECT 3.935 1.615 4.185 2.125 ;
        RECT 4.775 1.615 5.025 2.125 ;
        RECT 5.615 1.615 5.865 2.125 ;
        RECT 6.455 1.615 6.705 2.125 ;
        RECT 3.935 1.445 7.275 1.615 ;
        RECT 6.710 0.905 7.275 1.445 ;
        RECT 0.535 0.725 7.275 0.905 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 3.895 0.255 4.225 0.725 ;
        RECT 4.735 0.255 5.065 0.725 ;
        RECT 5.575 0.255 5.905 0.725 ;
        RECT 6.415 0.255 6.745 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.090 1.665 0.405 2.465 ;
        RECT 0.575 1.835 0.825 2.635 ;
        RECT 0.995 1.665 1.245 2.465 ;
        RECT 1.415 1.835 1.665 2.635 ;
        RECT 1.835 1.665 2.085 2.465 ;
        RECT 2.255 1.835 2.505 2.635 ;
        RECT 2.675 1.665 2.925 2.465 ;
        RECT 3.095 1.835 3.345 2.635 ;
        RECT 3.515 2.295 7.125 2.465 ;
        RECT 3.515 1.665 3.765 2.295 ;
        RECT 4.355 1.785 4.605 2.295 ;
        RECT 5.195 1.785 5.445 2.295 ;
        RECT 6.035 1.785 6.285 2.295 ;
        RECT 6.875 1.785 7.125 2.295 ;
        RECT 0.090 1.455 3.765 1.665 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.555 ;
        RECT 2.715 0.085 2.885 0.555 ;
        RECT 3.555 0.085 3.725 0.555 ;
        RECT 4.395 0.085 4.565 0.555 ;
        RECT 5.235 0.085 5.405 0.555 ;
        RECT 6.075 0.085 6.245 0.555 ;
        RECT 6.915 0.085 7.205 0.555 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
END sky130_fd_sc_hd__nor2_8

#--------EOF---------

MACRO sky130_fd_sc_hd__nor2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.960 1.065 1.325 1.325 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 0.725 0.325 1.325 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.725 0.785 2.075 1.015 ;
        RECT 0.240 0.105 2.075 0.785 ;
        RECT 0.240 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.435500 ;
    PORT
      LAYER li1 ;
        RECT 1.655 1.850 2.215 2.465 ;
        RECT 2.035 0.895 2.215 1.850 ;
        RECT 1.235 0.725 2.215 0.895 ;
        RECT 1.235 0.255 1.565 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.415 1.680 0.675 1.905 ;
        RECT 0.875 1.855 1.205 2.635 ;
        RECT 0.415 1.510 1.705 1.680 ;
        RECT 0.495 0.545 0.675 1.510 ;
        RECT 1.535 1.245 1.705 1.510 ;
        RECT 1.535 1.075 1.865 1.245 ;
        RECT 0.330 0.370 0.675 0.545 ;
        RECT 0.855 0.085 1.065 0.895 ;
        RECT 1.735 0.085 2.120 0.555 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__nor2b_1

#--------EOF---------

MACRO sky130_fd_sc_hd__nor2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.480 1.065 0.920 1.275 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.910 1.275 3.125 1.965 ;
        RECT 2.600 1.065 3.125 1.275 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.335 3.155 1.015 ;
        RECT 0.010 0.105 2.215 0.335 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.621000 ;
    PORT
      LAYER li1 ;
        RECT 1.415 0.895 1.665 2.125 ;
        RECT 0.535 0.725 1.705 0.895 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 1.375 0.255 1.705 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.655 0.405 2.465 ;
        RECT 0.575 1.825 0.825 2.635 ;
        RECT 0.995 2.295 2.125 2.465 ;
        RECT 0.995 1.655 1.245 2.295 ;
        RECT 0.085 1.445 1.245 1.655 ;
        RECT 1.835 1.890 2.125 2.295 ;
        RECT 1.835 1.445 2.090 1.890 ;
        RECT 2.395 1.615 2.565 2.460 ;
        RECT 2.775 2.145 3.025 2.635 ;
        RECT 2.260 1.445 2.565 1.615 ;
        RECT 2.260 1.245 2.430 1.445 ;
        RECT 1.875 1.075 2.430 1.245 ;
        RECT 2.215 0.895 2.430 1.075 ;
        RECT 0.085 0.085 0.365 0.895 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.895 ;
        RECT 2.215 0.725 2.565 0.895 ;
        RECT 2.395 0.445 2.565 0.725 ;
        RECT 2.775 0.085 3.030 0.845 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__nor2b_2

#--------EOF---------

MACRO sky130_fd_sc_hd__nor2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor2b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.360 1.075 1.800 1.275 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 4.445 1.075 4.975 1.320 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.875 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.242000 ;
    PORT
      LAYER li1 ;
        RECT 2.295 1.745 2.465 2.125 ;
        RECT 3.135 1.745 3.305 2.125 ;
        RECT 2.295 1.445 3.305 1.745 ;
        RECT 2.295 0.905 2.625 1.445 ;
        RECT 0.535 0.725 3.385 0.905 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 3.055 0.255 3.385 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.085 1.665 0.365 2.465 ;
        RECT 0.535 1.835 0.865 2.635 ;
        RECT 1.035 1.665 1.205 2.465 ;
        RECT 1.375 1.835 1.625 2.635 ;
        RECT 1.795 2.295 3.855 2.465 ;
        RECT 1.795 1.665 2.125 2.295 ;
        RECT 2.635 1.935 2.965 2.295 ;
        RECT 0.085 1.455 2.125 1.665 ;
        RECT 3.475 1.575 3.855 2.295 ;
        RECT 4.025 1.575 4.355 2.465 ;
        RECT 4.025 1.275 4.275 1.575 ;
        RECT 4.525 1.495 4.930 2.635 ;
        RECT 2.795 1.075 4.275 1.275 ;
        RECT 0.085 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.555 ;
        RECT 2.715 0.085 2.885 0.555 ;
        RECT 3.555 0.085 3.845 0.905 ;
        RECT 4.025 0.815 4.275 1.075 ;
        RECT 4.025 0.255 4.355 0.815 ;
        RECT 4.525 0.085 4.815 0.905 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
END sky130_fd_sc_hd__nor2b_4

#--------EOF---------

MACRO sky130_fd_sc_hd__nor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.485 0.655 1.755 1.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.325 0.830 2.005 ;
        RECT 0.595 0.995 0.975 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.995 0.425 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.775 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.604500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 2.280 1.170 2.450 ;
        RECT 0.090 1.495 0.425 2.280 ;
        RECT 1.000 1.665 1.170 2.280 ;
        RECT 1.000 1.495 1.315 1.665 ;
        RECT 1.145 0.825 1.315 1.495 ;
        RECT 0.090 0.655 1.315 0.825 ;
        RECT 0.090 0.385 0.345 0.655 ;
        RECT 1.015 0.385 1.185 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 1.435 1.835 1.750 2.635 ;
        RECT 0.515 0.085 0.845 0.485 ;
        RECT 1.355 0.085 1.685 0.485 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__nor3_1

#--------EOF---------

MACRO sky130_fd_sc_hd__nor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.135 1.075 0.965 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.135 1.075 2.185 1.285 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.375 1.285 2.640 1.625 ;
        RECT 2.375 1.075 2.965 1.285 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.105 3.595 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.796500 ;
    PORT
      LAYER li1 ;
        RECT 2.835 1.625 3.045 2.125 ;
        RECT 2.835 1.455 3.595 1.625 ;
        RECT 3.135 0.905 3.595 1.455 ;
        RECT 0.535 0.725 3.595 0.905 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.755 0.255 3.085 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.150 1.625 0.405 2.465 ;
        RECT 0.575 1.795 0.825 2.635 ;
        RECT 0.995 1.625 1.245 2.465 ;
        RECT 1.415 2.295 3.465 2.465 ;
        RECT 1.415 1.795 1.665 2.295 ;
        RECT 1.835 1.625 2.085 2.125 ;
        RECT 2.415 1.795 2.625 2.295 ;
        RECT 3.215 1.795 3.465 2.295 ;
        RECT 0.150 1.455 2.085 1.625 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.585 0.555 ;
        RECT 3.255 0.085 3.545 0.555 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__nor3_2

#--------EOF---------

MACRO sky130_fd_sc_hd__nor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 1.825 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.515 1.445 5.165 1.615 ;
        RECT 3.515 1.285 3.685 1.445 ;
        RECT 2.095 1.075 3.685 1.285 ;
        RECT 4.995 1.285 5.165 1.445 ;
        RECT 4.995 1.075 5.415 1.285 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.855 1.075 4.765 1.275 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.575 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.593000 ;
    PORT
      LAYER li1 ;
        RECT 3.515 1.965 3.765 2.125 ;
        RECT 4.355 1.965 4.605 2.125 ;
        RECT 3.515 1.955 4.605 1.965 ;
        RECT 5.615 1.955 5.895 2.465 ;
        RECT 3.515 1.785 5.895 1.955 ;
        RECT 5.605 0.905 5.895 1.785 ;
        RECT 0.535 0.725 5.895 0.905 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 3.895 0.255 4.225 0.725 ;
        RECT 4.735 0.255 5.065 0.725 ;
        RECT 5.605 0.255 5.895 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.150 1.625 0.405 2.465 ;
        RECT 0.575 1.795 0.825 2.635 ;
        RECT 0.995 1.625 1.245 2.465 ;
        RECT 1.415 1.795 1.665 2.635 ;
        RECT 1.835 2.085 2.925 2.465 ;
        RECT 1.835 1.625 2.085 2.085 ;
        RECT 0.150 1.455 2.085 1.625 ;
        RECT 2.255 1.625 2.505 1.915 ;
        RECT 2.675 1.795 2.925 2.085 ;
        RECT 3.095 2.295 5.025 2.465 ;
        RECT 3.095 1.625 3.345 2.295 ;
        RECT 3.935 2.135 4.185 2.295 ;
        RECT 4.775 2.135 5.025 2.295 ;
        RECT 5.195 2.125 5.445 2.465 ;
        RECT 2.255 1.455 3.345 1.625 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.555 ;
        RECT 2.715 0.085 2.885 0.555 ;
        RECT 3.555 0.085 3.725 0.555 ;
        RECT 4.395 0.085 4.565 0.555 ;
        RECT 5.235 0.085 5.405 0.555 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 2.445 2.125 2.615 2.295 ;
        RECT 5.205 2.125 5.375 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
      LAYER met1 ;
        RECT 2.385 2.280 2.680 2.335 ;
        RECT 5.145 2.280 5.440 2.335 ;
        RECT 2.385 2.140 5.440 2.280 ;
        RECT 2.385 2.065 2.680 2.140 ;
        RECT 5.145 2.065 5.440 2.140 ;
  END
END sky130_fd_sc_hd__nor3_4

#--------EOF---------

MACRO sky130_fd_sc_hd__nor3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.475 0.995 1.815 1.615 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.065 0.995 1.305 1.615 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.995 2.335 1.615 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.185 0.335 2.520 1.015 ;
        RECT 0.185 0.105 2.035 0.335 ;
        RECT 0.185 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.716500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.445 0.545 2.455 ;
        RECT 0.085 0.825 0.255 1.445 ;
        RECT 0.085 0.655 1.445 0.825 ;
        RECT 0.085 0.255 0.605 0.655 ;
        RECT 1.275 0.310 1.445 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 1.615 2.125 1.945 2.635 ;
        RECT 0.715 1.785 2.675 1.955 ;
        RECT 0.715 1.245 0.885 1.785 ;
        RECT 0.425 1.075 0.885 1.245 ;
        RECT 2.505 0.825 2.675 1.785 ;
        RECT 0.775 0.085 1.105 0.485 ;
        RECT 1.615 0.085 1.945 0.825 ;
        RECT 2.180 0.655 2.675 0.825 ;
        RECT 2.180 0.405 2.350 0.655 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__nor3b_1

#--------EOF---------

MACRO sky130_fd_sc_hd__nor3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.965 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.135 1.075 2.640 1.285 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 4.030 1.075 4.515 1.285 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 4.595 1.015 ;
        RECT 0.005 0.105 3.635 0.335 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.796500 ;
    PORT
      LAYER li1 ;
        RECT 2.815 0.905 3.065 2.125 ;
        RECT 0.535 0.725 3.105 0.905 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.775 0.255 3.105 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.090 1.625 0.405 2.465 ;
        RECT 0.575 1.795 0.825 2.635 ;
        RECT 0.995 1.625 1.245 2.465 ;
        RECT 1.415 2.295 3.480 2.465 ;
        RECT 1.415 1.795 1.665 2.295 ;
        RECT 1.835 1.625 2.085 2.125 ;
        RECT 0.090 1.455 2.085 1.625 ;
        RECT 2.375 1.455 2.645 2.295 ;
        RECT 3.235 1.455 3.480 2.295 ;
        RECT 3.690 1.455 4.045 1.870 ;
        RECT 4.215 1.540 4.465 2.635 ;
        RECT 3.690 1.285 3.860 1.455 ;
        RECT 3.235 1.075 3.860 1.285 ;
        RECT 3.690 0.905 3.860 1.075 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.605 0.555 ;
        RECT 3.275 0.085 3.480 0.895 ;
        RECT 3.690 0.380 4.045 0.905 ;
        RECT 4.215 0.085 4.505 0.825 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__nor3b_2

#--------EOF---------

MACRO sky130_fd_sc_hd__nor3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor3b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.035 1.075 2.690 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.035 1.075 4.300 1.285 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.445 1.285 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.515 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.593000 ;
    PORT
      LAYER li1 ;
        RECT 4.875 1.625 5.125 2.125 ;
        RECT 5.715 1.625 5.965 2.125 ;
        RECT 6.555 1.625 6.760 2.415 ;
        RECT 4.875 1.455 6.760 1.625 ;
        RECT 6.420 0.905 6.760 1.455 ;
        RECT 0.955 0.725 6.760 0.905 ;
        RECT 0.955 0.255 1.285 0.725 ;
        RECT 1.795 0.255 2.125 0.725 ;
        RECT 3.155 0.255 3.485 0.725 ;
        RECT 3.995 0.255 4.325 0.725 ;
        RECT 4.835 0.255 5.165 0.725 ;
        RECT 5.675 0.255 6.005 0.725 ;
        RECT 6.515 0.315 6.760 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.110 1.625 0.405 2.465 ;
        RECT 0.575 1.795 0.825 2.635 ;
        RECT 0.995 1.965 1.245 2.465 ;
        RECT 1.415 2.135 1.665 2.635 ;
        RECT 1.835 1.965 2.085 2.465 ;
        RECT 2.255 2.135 2.505 2.635 ;
        RECT 2.775 2.295 6.385 2.465 ;
        RECT 2.775 2.135 3.025 2.295 ;
        RECT 3.615 2.135 3.865 2.295 ;
        RECT 3.195 1.965 3.445 2.125 ;
        RECT 4.035 1.965 4.285 2.125 ;
        RECT 0.995 1.795 4.285 1.965 ;
        RECT 4.455 1.795 4.705 2.295 ;
        RECT 5.295 1.795 5.545 2.295 ;
        RECT 6.135 1.795 6.385 2.295 ;
        RECT 0.110 1.455 4.705 1.625 ;
        RECT 0.615 0.905 0.785 1.455 ;
        RECT 4.535 1.285 4.705 1.455 ;
        RECT 4.535 1.075 6.125 1.285 ;
        RECT 0.110 0.735 0.785 0.905 ;
        RECT 0.110 0.255 0.445 0.735 ;
        RECT 0.615 0.085 0.785 0.555 ;
        RECT 1.455 0.085 1.625 0.555 ;
        RECT 2.295 0.085 2.985 0.555 ;
        RECT 3.655 0.085 3.825 0.555 ;
        RECT 4.495 0.085 4.665 0.555 ;
        RECT 5.335 0.085 5.505 0.555 ;
        RECT 6.175 0.085 6.345 0.555 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
  END
END sky130_fd_sc_hd__nor3b_4

#--------EOF---------

MACRO sky130_fd_sc_hd__nor4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.955 0.655 2.215 1.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.455 1.245 1.695 2.450 ;
        RECT 1.245 1.075 1.695 1.245 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.030 1.615 1.285 2.450 ;
        RECT 0.845 1.415 1.285 1.615 ;
        RECT 0.845 0.995 1.075 1.415 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.745 0.335 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.295 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.672750 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.665 0.425 2.450 ;
        RECT 0.090 1.495 0.675 1.665 ;
        RECT 0.505 0.825 0.675 1.495 ;
        RECT 0.505 0.655 1.705 0.825 ;
        RECT 0.505 0.645 0.860 0.655 ;
        RECT 0.595 0.385 0.860 0.645 ;
        RECT 1.535 0.385 1.705 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 1.955 1.835 2.215 2.635 ;
        RECT 0.085 0.085 0.345 0.575 ;
        RECT 1.035 0.085 1.365 0.485 ;
        RECT 1.875 0.085 2.205 0.485 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__nor4_1

#--------EOF---------

MACRO sky130_fd_sc_hd__nor4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.200 1.075 0.965 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.135 1.075 1.940 1.285 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.210 1.075 3.105 1.285 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.340 1.075 3.925 1.285 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.455 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.972000 ;
    PORT
      LAYER li1 ;
        RECT 3.655 1.625 3.905 2.125 ;
        RECT 3.655 1.455 4.515 1.625 ;
        RECT 4.180 0.905 4.515 1.455 ;
        RECT 0.535 0.725 4.515 0.905 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.775 0.255 3.105 0.725 ;
        RECT 3.615 0.255 3.945 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.150 1.625 0.405 2.465 ;
        RECT 0.575 1.795 0.825 2.635 ;
        RECT 0.995 1.625 1.245 2.465 ;
        RECT 1.415 2.295 3.065 2.465 ;
        RECT 1.415 1.795 1.665 2.295 ;
        RECT 1.835 1.625 2.085 2.125 ;
        RECT 0.150 1.455 2.085 1.625 ;
        RECT 2.395 1.625 2.645 2.125 ;
        RECT 2.815 1.795 3.065 2.295 ;
        RECT 3.235 2.295 4.325 2.465 ;
        RECT 3.235 1.625 3.485 2.295 ;
        RECT 4.075 1.795 4.325 2.295 ;
        RECT 2.395 1.455 3.485 1.625 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.605 0.555 ;
        RECT 3.275 0.085 3.445 0.555 ;
        RECT 4.115 0.085 4.405 0.555 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__nor4_2

#--------EOF---------

MACRO sky130_fd_sc_hd__nor4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.180 1.075 1.825 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 2.095 1.075 4.070 1.285 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 4.295 1.075 5.705 1.285 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 5.875 1.075 7.295 1.285 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.775 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.944000 ;
    PORT
      LAYER li1 ;
        RECT 6.135 1.625 6.385 2.125 ;
        RECT 6.975 1.625 7.225 2.125 ;
        RECT 6.135 1.455 7.735 1.625 ;
        RECT 7.465 0.905 7.735 1.455 ;
        RECT 0.535 0.725 7.735 0.905 ;
        RECT 0.535 0.255 0.865 0.725 ;
        RECT 1.375 0.255 1.705 0.725 ;
        RECT 2.215 0.255 2.545 0.725 ;
        RECT 3.055 0.255 3.385 0.725 ;
        RECT 4.415 0.255 4.745 0.725 ;
        RECT 5.255 0.255 5.585 0.725 ;
        RECT 6.095 0.255 6.425 0.725 ;
        RECT 6.935 0.255 7.265 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.090 1.625 0.405 2.465 ;
        RECT 0.575 1.795 0.825 2.635 ;
        RECT 0.995 1.625 1.245 2.465 ;
        RECT 1.415 1.795 1.665 2.635 ;
        RECT 1.835 2.295 3.820 2.465 ;
        RECT 1.835 1.625 2.085 2.295 ;
        RECT 0.090 1.455 2.085 1.625 ;
        RECT 2.255 1.625 2.505 2.125 ;
        RECT 2.675 1.795 2.925 2.295 ;
        RECT 3.095 1.625 3.345 2.125 ;
        RECT 3.515 1.795 3.820 2.295 ;
        RECT 4.005 2.295 7.645 2.465 ;
        RECT 4.005 1.795 4.285 2.295 ;
        RECT 4.455 1.625 4.705 2.125 ;
        RECT 4.875 1.795 5.125 2.295 ;
        RECT 5.295 1.625 5.545 2.125 ;
        RECT 5.715 1.795 5.965 2.295 ;
        RECT 6.555 1.795 6.805 2.295 ;
        RECT 7.395 1.795 7.645 2.295 ;
        RECT 2.255 1.455 5.545 1.625 ;
        RECT 0.090 0.085 0.365 0.905 ;
        RECT 1.035 0.085 1.205 0.555 ;
        RECT 1.875 0.085 2.045 0.555 ;
        RECT 2.715 0.085 2.885 0.555 ;
        RECT 3.555 0.085 4.245 0.555 ;
        RECT 4.915 0.085 5.085 0.555 ;
        RECT 5.755 0.085 5.925 0.555 ;
        RECT 6.595 0.085 6.765 0.555 ;
        RECT 7.435 0.085 7.605 0.555 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
  END
END sky130_fd_sc_hd__nor4_4

#--------EOF---------

MACRO sky130_fd_sc_hd__nor4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.955 0.995 2.275 1.615 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.455 0.995 1.785 1.615 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.985 0.995 1.285 1.615 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.995 2.795 1.615 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.245 0.335 3.000 1.015 ;
        RECT 0.245 0.105 2.515 0.335 ;
        RECT 0.245 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.871000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.825 0.345 2.450 ;
        RECT 0.085 0.655 1.925 0.825 ;
        RECT 0.855 0.300 1.055 0.655 ;
        RECT 1.725 0.310 1.925 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 2.095 2.185 2.425 2.635 ;
        RECT 0.525 1.795 3.135 2.005 ;
        RECT 0.525 0.995 0.745 1.795 ;
        RECT 2.965 0.825 3.135 1.795 ;
        RECT 0.355 0.085 0.685 0.480 ;
        RECT 1.225 0.085 1.555 0.485 ;
        RECT 2.095 0.085 2.425 0.825 ;
        RECT 2.660 0.655 3.135 0.825 ;
        RECT 2.660 0.405 2.830 0.655 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__nor4b_1

#--------EOF---------

MACRO sky130_fd_sc_hd__nor4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.100 1.075 1.240 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.420 1.075 2.635 1.285 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.815 1.075 3.535 1.285 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 5.185 1.285 5.435 1.955 ;
        RECT 4.805 1.075 5.435 1.285 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 5.370 1.015 ;
        RECT 0.005 0.105 4.430 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.972000 ;
    PORT
      LAYER li1 ;
        RECT 3.630 1.625 3.880 2.125 ;
        RECT 3.630 1.455 4.035 1.625 ;
        RECT 3.715 1.075 4.035 1.455 ;
        RECT 3.715 0.905 3.920 1.075 ;
        RECT 0.515 0.725 3.920 0.905 ;
        RECT 0.515 0.255 0.845 0.725 ;
        RECT 1.355 0.255 1.685 0.725 ;
        RECT 2.750 0.255 3.080 0.725 ;
        RECT 3.590 0.255 3.920 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.085 1.625 0.425 2.465 ;
        RECT 0.595 1.795 0.805 2.635 ;
        RECT 0.975 1.625 1.225 2.465 ;
        RECT 1.395 2.295 3.040 2.465 ;
        RECT 1.395 1.795 1.605 2.295 ;
        RECT 1.775 1.625 2.105 2.125 ;
        RECT 0.085 1.455 2.105 1.625 ;
        RECT 2.275 1.625 2.660 2.125 ;
        RECT 2.830 1.795 3.040 2.295 ;
        RECT 3.210 2.295 4.295 2.465 ;
        RECT 3.210 1.625 3.460 2.295 ;
        RECT 4.050 1.795 4.295 2.295 ;
        RECT 4.465 2.035 4.820 2.450 ;
        RECT 4.990 2.135 5.240 2.635 ;
        RECT 2.275 1.455 3.460 1.625 ;
        RECT 4.465 1.245 4.635 2.035 ;
        RECT 4.320 1.075 4.635 1.245 ;
        RECT 4.465 0.905 4.635 1.075 ;
        RECT 0.085 0.085 0.345 0.905 ;
        RECT 1.015 0.085 1.185 0.555 ;
        RECT 1.855 0.085 2.580 0.555 ;
        RECT 3.250 0.085 3.420 0.555 ;
        RECT 4.090 0.085 4.295 0.895 ;
        RECT 4.465 0.380 4.820 0.905 ;
        RECT 4.990 0.085 5.240 0.825 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__nor4b_2

#--------EOF---------

MACRO sky130_fd_sc_hd__nor4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.395 1.075 1.805 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 2.075 1.075 3.750 1.285 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.985 1.075 5.685 1.285 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 7.810 1.075 8.655 1.285 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 8.715 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.944000 ;
    PORT
      LAYER li1 ;
        RECT 6.115 1.625 6.365 2.125 ;
        RECT 6.955 1.625 7.205 2.125 ;
        RECT 6.115 1.455 7.205 1.625 ;
        RECT 6.115 0.905 6.465 1.455 ;
        RECT 0.515 0.725 7.245 0.905 ;
        RECT 0.515 0.255 0.845 0.725 ;
        RECT 1.355 0.255 1.685 0.725 ;
        RECT 2.195 0.255 2.525 0.725 ;
        RECT 3.035 0.255 3.365 0.725 ;
        RECT 4.395 0.255 4.725 0.725 ;
        RECT 5.235 0.255 5.565 0.725 ;
        RECT 6.075 0.255 6.405 0.725 ;
        RECT 6.915 0.255 7.245 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.740 2.805 ;
        RECT 0.095 1.625 0.425 2.465 ;
        RECT 0.595 1.795 0.805 2.635 ;
        RECT 0.975 1.625 1.225 2.465 ;
        RECT 1.395 1.795 1.645 2.635 ;
        RECT 1.815 2.295 3.745 2.465 ;
        RECT 1.815 1.625 2.065 2.295 ;
        RECT 0.095 1.455 2.065 1.625 ;
        RECT 2.235 1.625 2.485 2.125 ;
        RECT 2.655 1.795 2.905 2.295 ;
        RECT 3.075 1.625 3.325 2.125 ;
        RECT 3.495 1.795 3.745 2.295 ;
        RECT 4.015 2.295 7.625 2.465 ;
        RECT 4.015 1.795 4.265 2.295 ;
        RECT 4.435 1.625 4.685 2.125 ;
        RECT 4.855 1.795 5.105 2.295 ;
        RECT 5.275 1.625 5.525 2.125 ;
        RECT 2.235 1.455 5.525 1.625 ;
        RECT 5.695 1.455 5.945 2.295 ;
        RECT 6.535 1.795 6.785 2.295 ;
        RECT 7.375 1.795 7.625 2.295 ;
        RECT 7.850 1.625 8.185 2.465 ;
        RECT 7.470 1.455 8.185 1.625 ;
        RECT 8.355 1.455 8.585 2.635 ;
        RECT 7.470 1.285 7.640 1.455 ;
        RECT 6.635 1.075 7.640 1.285 ;
        RECT 7.470 0.905 7.640 1.075 ;
        RECT 0.175 0.085 0.345 0.895 ;
        RECT 7.470 0.735 8.185 0.905 ;
        RECT 1.015 0.085 1.185 0.555 ;
        RECT 1.855 0.085 2.025 0.555 ;
        RECT 2.695 0.085 2.865 0.555 ;
        RECT 3.535 0.085 4.225 0.555 ;
        RECT 4.895 0.085 5.065 0.555 ;
        RECT 5.735 0.085 5.905 0.555 ;
        RECT 6.575 0.085 6.745 0.555 ;
        RECT 7.415 0.085 7.585 0.555 ;
        RECT 7.810 0.255 8.185 0.735 ;
        RECT 8.355 0.085 8.585 0.905 ;
        RECT 0.000 -0.085 8.740 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
  END
END sky130_fd_sc_hd__nor4b_4

#--------EOF---------

MACRO sky130_fd_sc_hd__nor4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4bb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.295 1.275 3.595 1.705 ;
        RECT 3.115 0.995 3.595 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.825 1.630 3.085 2.410 ;
        RECT 2.615 1.445 3.085 1.630 ;
        RECT 2.615 0.995 2.945 1.445 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.430 0.995 0.780 1.695 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.950 0.995 1.240 1.325 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.045 0.335 3.675 1.015 ;
        RECT 0.150 -0.085 0.320 0.335 ;
        RECT 1.425 0.105 3.675 0.335 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.606900 ;
    PORT
      LAYER li1 ;
        RECT 1.470 1.955 2.055 2.125 ;
        RECT 1.855 0.825 2.055 1.955 ;
        RECT 1.855 0.655 3.085 0.825 ;
        RECT 2.015 0.300 2.215 0.655 ;
        RECT 2.885 0.310 3.085 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 2.070 0.345 2.455 ;
        RECT 0.515 2.240 0.845 2.635 ;
        RECT 1.035 2.295 2.395 2.465 ;
        RECT 1.035 2.070 1.205 2.295 ;
        RECT 0.085 1.885 1.205 2.070 ;
        RECT 0.085 0.825 0.260 1.885 ;
        RECT 0.995 1.525 1.590 1.715 ;
        RECT 1.410 1.325 1.590 1.525 ;
        RECT 1.410 0.995 1.685 1.325 ;
        RECT 2.225 0.995 2.395 2.295 ;
        RECT 3.255 1.875 3.585 2.635 ;
        RECT 1.410 0.825 1.590 0.995 ;
        RECT 0.085 0.450 0.405 0.825 ;
        RECT 0.655 0.085 0.825 0.825 ;
        RECT 1.075 0.655 1.590 0.825 ;
        RECT 1.075 0.450 1.245 0.655 ;
        RECT 1.515 0.085 1.845 0.480 ;
        RECT 2.385 0.085 2.715 0.485 ;
        RECT 3.255 0.085 3.585 0.825 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__nor4bb_1

#--------EOF---------

MACRO sky130_fd_sc_hd__nor4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4bb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 5.130 1.075 5.895 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.165 1.075 4.960 1.275 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.950 0.995 1.235 1.325 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.780 1.695 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.045 0.335 5.975 1.015 ;
        RECT 0.145 -0.085 0.315 0.335 ;
        RECT 1.470 0.105 5.975 0.335 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.972000 ;
    PORT
      LAYER li1 ;
        RECT 2.900 1.445 3.995 1.705 ;
        RECT 3.575 0.905 3.995 1.445 ;
        RECT 2.060 0.725 5.450 0.905 ;
        RECT 2.060 0.255 2.390 0.725 ;
        RECT 2.900 0.255 3.230 0.725 ;
        RECT 4.280 0.255 4.610 0.725 ;
        RECT 5.120 0.255 5.450 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.085 2.055 0.345 2.455 ;
        RECT 0.515 2.240 0.845 2.635 ;
        RECT 1.640 2.295 3.650 2.465 ;
        RECT 1.640 2.225 1.970 2.295 ;
        RECT 2.480 2.215 3.650 2.295 ;
        RECT 3.860 2.215 4.990 2.465 ;
        RECT 0.085 1.885 1.915 2.055 ;
        RECT 0.085 0.825 0.255 1.885 ;
        RECT 0.995 1.525 1.575 1.715 ;
        RECT 1.405 1.245 1.575 1.525 ;
        RECT 1.745 1.585 1.915 1.885 ;
        RECT 2.140 2.045 2.310 2.125 ;
        RECT 2.140 1.875 4.610 2.045 ;
        RECT 2.140 1.795 2.310 1.875 ;
        RECT 1.745 1.415 2.730 1.585 ;
        RECT 4.320 1.455 4.610 1.875 ;
        RECT 4.780 1.625 4.990 2.215 ;
        RECT 5.160 1.795 5.370 2.635 ;
        RECT 5.540 1.625 5.870 2.465 ;
        RECT 4.780 1.455 5.870 1.625 ;
        RECT 2.560 1.275 2.730 1.415 ;
        RECT 1.405 1.075 2.390 1.245 ;
        RECT 2.560 1.075 3.405 1.275 ;
        RECT 1.405 0.825 1.575 1.075 ;
        RECT 0.085 0.450 0.465 0.825 ;
        RECT 0.635 0.085 0.805 0.825 ;
        RECT 1.055 0.655 1.575 0.825 ;
        RECT 1.055 0.450 1.250 0.655 ;
        RECT 1.560 0.085 1.890 0.480 ;
        RECT 2.560 0.085 2.730 0.555 ;
        RECT 3.400 0.085 4.110 0.555 ;
        RECT 4.780 0.085 4.950 0.555 ;
        RECT 5.620 0.085 5.895 0.905 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
END sky130_fd_sc_hd__nor4bb_2

#--------EOF---------

MACRO sky130_fd_sc_hd__nor4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__nor4bb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 7.375 1.075 9.110 1.285 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 5.150 1.075 7.105 1.285 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 0.445 1.365 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.955 1.075 1.295 1.325 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.105 9.195 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.390 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.944000 ;
    PORT
      LAYER li1 ;
        RECT 1.840 1.415 3.185 1.705 ;
        RECT 3.015 0.905 3.185 1.415 ;
        RECT 1.935 0.725 8.665 0.905 ;
        RECT 1.935 0.255 2.265 0.725 ;
        RECT 2.775 0.255 3.105 0.725 ;
        RECT 3.615 0.255 3.945 0.725 ;
        RECT 4.455 0.255 4.785 0.725 ;
        RECT 5.815 0.255 6.145 0.725 ;
        RECT 6.655 0.255 6.985 0.725 ;
        RECT 7.495 0.255 7.825 0.725 ;
        RECT 8.335 0.255 8.665 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.085 2.045 0.365 2.465 ;
        RECT 0.535 2.215 0.865 2.635 ;
        RECT 1.515 2.295 5.195 2.465 ;
        RECT 1.515 2.215 3.525 2.295 ;
        RECT 0.085 1.875 3.525 2.045 ;
        RECT 0.085 1.535 0.785 1.875 ;
        RECT 0.955 1.535 1.635 1.705 ;
        RECT 0.615 0.895 0.785 1.535 ;
        RECT 1.465 1.245 1.635 1.535 ;
        RECT 3.355 1.285 3.525 1.875 ;
        RECT 3.695 1.625 3.905 2.125 ;
        RECT 4.075 1.795 4.325 2.295 ;
        RECT 4.495 1.625 4.745 2.125 ;
        RECT 4.915 1.795 5.195 2.295 ;
        RECT 5.380 2.295 7.365 2.465 ;
        RECT 5.380 1.795 5.685 2.295 ;
        RECT 5.855 1.625 6.105 2.125 ;
        RECT 6.275 1.795 6.525 2.295 ;
        RECT 6.695 1.625 6.945 2.125 ;
        RECT 3.695 1.455 6.945 1.625 ;
        RECT 7.115 1.625 7.365 2.295 ;
        RECT 7.535 1.795 7.785 2.635 ;
        RECT 7.955 1.625 8.205 2.465 ;
        RECT 8.375 1.795 8.625 2.635 ;
        RECT 8.795 1.625 9.110 2.465 ;
        RECT 7.115 1.455 9.110 1.625 ;
        RECT 1.465 1.075 2.845 1.245 ;
        RECT 3.355 1.075 4.905 1.285 ;
        RECT 1.465 0.905 1.635 1.075 ;
        RECT 0.085 0.725 0.785 0.895 ;
        RECT 0.955 0.735 1.635 0.905 ;
        RECT 0.085 0.255 0.445 0.725 ;
        RECT 0.615 0.085 0.785 0.555 ;
        RECT 0.955 0.255 1.285 0.735 ;
        RECT 1.595 0.085 1.765 0.555 ;
        RECT 2.435 0.085 2.605 0.555 ;
        RECT 3.275 0.085 3.445 0.555 ;
        RECT 4.115 0.085 4.285 0.555 ;
        RECT 4.955 0.085 5.645 0.555 ;
        RECT 6.315 0.085 6.485 0.555 ;
        RECT 7.155 0.085 7.325 0.555 ;
        RECT 7.995 0.085 8.165 0.555 ;
        RECT 8.835 0.085 9.110 0.905 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
  END
END sky130_fd_sc_hd__nor4bb_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o2bb2a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.770 1.075 1.220 1.275 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.390 0.905 1.565 1.100 ;
        RECT 1.070 0.735 1.565 0.905 ;
        RECT 1.070 0.380 1.290 0.735 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 3.250 1.075 3.595 1.645 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.325 3.080 2.425 ;
        RECT 2.520 1.075 3.080 1.325 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 0.930 1.015 ;
        RECT 0.005 0.105 3.675 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.795 0.345 2.465 ;
        RECT 0.085 0.825 0.260 1.795 ;
        RECT 0.085 0.255 0.425 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.515 2.235 0.845 2.635 ;
        RECT 1.715 2.235 2.115 2.635 ;
        RECT 2.405 2.055 2.735 2.290 ;
        RECT 0.655 1.885 2.735 2.055 ;
        RECT 0.655 1.615 0.825 1.885 ;
        RECT 0.430 1.445 0.825 1.615 ;
        RECT 0.995 1.495 2.010 1.715 ;
        RECT 0.430 0.995 0.600 1.445 ;
        RECT 1.735 1.355 2.010 1.495 ;
        RECT 2.180 1.495 2.735 1.885 ;
        RECT 3.250 1.815 3.595 2.635 ;
        RECT 0.620 0.085 0.790 0.750 ;
        RECT 1.735 0.565 1.905 1.355 ;
        RECT 2.180 1.245 2.350 1.495 ;
        RECT 2.155 1.075 2.350 1.245 ;
        RECT 2.155 0.690 2.325 1.075 ;
        RECT 1.460 0.395 1.905 0.565 ;
        RECT 2.075 0.320 2.325 0.690 ;
        RECT 2.495 0.725 3.595 0.905 ;
        RECT 2.495 0.320 2.745 0.725 ;
        RECT 2.915 0.085 3.085 0.555 ;
        RECT 3.255 0.320 3.595 0.725 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__o2bb2a_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o2bb2a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.215 1.075 1.685 1.275 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.855 0.905 2.025 1.100 ;
        RECT 1.515 0.770 2.025 0.905 ;
        RECT 1.515 0.735 2.020 0.770 ;
        RECT 1.515 0.380 1.735 0.735 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 3.700 1.075 4.045 1.645 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 3.355 1.325 3.525 2.425 ;
        RECT 2.970 1.075 3.525 1.325 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.785 1.375 1.015 ;
        RECT 0.005 0.105 4.135 0.785 ;
        RECT 0.135 -0.085 0.305 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.535 1.795 0.790 2.465 ;
        RECT 0.535 0.825 0.705 1.795 ;
        RECT 0.535 0.255 0.870 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.110 1.410 0.365 2.635 ;
        RECT 0.960 2.235 1.290 2.635 ;
        RECT 2.160 2.235 2.565 2.635 ;
        RECT 2.835 2.055 3.185 2.425 ;
        RECT 1.100 1.885 3.185 2.055 ;
        RECT 1.100 1.615 1.270 1.885 ;
        RECT 0.875 1.445 1.270 1.615 ;
        RECT 1.440 1.495 2.460 1.715 ;
        RECT 0.875 0.995 1.045 1.445 ;
        RECT 2.195 1.355 2.460 1.495 ;
        RECT 2.630 1.495 3.185 1.885 ;
        RECT 3.730 1.815 4.045 2.635 ;
        RECT 0.110 0.085 0.365 0.910 ;
        RECT 1.065 0.085 1.235 0.750 ;
        RECT 2.195 0.565 2.365 1.355 ;
        RECT 2.630 1.245 2.800 1.495 ;
        RECT 2.610 1.075 2.800 1.245 ;
        RECT 2.610 0.690 2.780 1.075 ;
        RECT 1.905 0.395 2.365 0.565 ;
        RECT 2.535 0.320 2.780 0.690 ;
        RECT 2.955 0.725 4.045 0.905 ;
        RECT 2.955 0.320 3.185 0.725 ;
        RECT 3.375 0.085 3.545 0.555 ;
        RECT 3.715 0.320 4.045 0.725 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__o2bb2a_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o2bb2a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.315 1.445 4.965 1.615 ;
        RECT 3.315 1.075 3.645 1.445 ;
        RECT 4.605 1.075 4.965 1.445 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.815 1.075 4.435 1.275 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.445 1.895 1.615 ;
        RECT 0.085 1.075 0.575 1.445 ;
        RECT 1.565 1.075 1.895 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.805 1.075 1.345 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.915 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 5.275 1.955 5.525 2.465 ;
        RECT 6.115 1.955 6.365 2.465 ;
        RECT 5.275 1.785 6.365 1.955 ;
        RECT 6.115 1.655 6.365 1.785 ;
        RECT 6.115 1.415 6.910 1.655 ;
        RECT 6.605 0.905 6.910 1.415 ;
        RECT 5.235 0.725 6.910 0.905 ;
        RECT 5.235 0.275 5.565 0.725 ;
        RECT 6.075 0.275 6.405 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.140 1.795 0.345 2.635 ;
        RECT 0.555 2.295 1.645 2.465 ;
        RECT 0.555 1.785 0.805 2.295 ;
        RECT 1.395 2.125 1.645 2.295 ;
        RECT 1.815 2.125 2.065 2.635 ;
        RECT 0.975 1.955 1.225 2.125 ;
        RECT 2.235 1.965 2.525 2.465 ;
        RECT 2.695 2.135 3.425 2.635 ;
        RECT 4.015 2.135 4.265 2.635 ;
        RECT 3.595 1.965 3.845 2.125 ;
        RECT 4.435 1.965 4.685 2.465 ;
        RECT 2.235 1.955 2.615 1.965 ;
        RECT 0.975 1.785 2.615 1.955 ;
        RECT 2.065 1.415 2.615 1.785 ;
        RECT 2.955 1.785 4.685 1.965 ;
        RECT 4.855 1.795 5.105 2.635 ;
        RECT 5.695 2.165 5.945 2.635 ;
        RECT 6.535 1.825 6.785 2.635 ;
        RECT 2.065 1.075 2.445 1.415 ;
        RECT 2.955 1.245 3.145 1.785 ;
        RECT 2.615 1.075 3.145 1.245 ;
        RECT 5.165 1.245 5.455 1.615 ;
        RECT 5.165 1.075 6.435 1.245 ;
        RECT 0.095 0.735 2.025 0.905 ;
        RECT 0.095 0.725 1.265 0.735 ;
        RECT 0.095 0.255 0.425 0.725 ;
        RECT 0.595 0.085 0.765 0.555 ;
        RECT 0.935 0.255 1.265 0.725 ;
        RECT 1.435 0.085 1.605 0.555 ;
        RECT 1.775 0.475 2.025 0.735 ;
        RECT 2.195 0.815 2.445 1.075 ;
        RECT 2.955 0.905 3.145 1.075 ;
        RECT 2.195 0.645 2.525 0.815 ;
        RECT 2.955 0.725 4.305 0.905 ;
        RECT 3.975 0.645 4.305 0.725 ;
        RECT 1.775 0.255 2.945 0.475 ;
        RECT 3.215 0.085 3.385 0.555 ;
        RECT 4.475 0.475 4.725 0.895 ;
        RECT 3.555 0.305 4.725 0.475 ;
        RECT 4.895 0.085 5.065 0.895 ;
        RECT 5.735 0.085 5.905 0.555 ;
        RECT 6.575 0.085 6.745 0.555 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 2.445 1.445 2.615 1.615 ;
        RECT 5.225 1.445 5.395 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
      LAYER met1 ;
        RECT 2.385 1.600 2.675 1.645 ;
        RECT 5.165 1.600 5.455 1.645 ;
        RECT 2.385 1.460 5.455 1.600 ;
        RECT 2.385 1.415 2.675 1.460 ;
        RECT 5.165 1.415 5.455 1.460 ;
  END
END sky130_fd_sc_hd__o2bb2a_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o2bb2ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.985 0.435 1.285 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 0.995 1.000 1.325 ;
        RECT 0.605 0.280 0.825 0.995 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.785 1.075 3.135 1.285 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.325 2.615 2.425 ;
        RECT 2.030 1.075 2.615 1.325 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.200 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 1.940 1.665 2.270 2.465 ;
        RECT 1.640 1.495 2.270 1.665 ;
        RECT 1.640 0.790 1.810 1.495 ;
        RECT 1.560 0.430 1.810 0.790 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.150 1.455 0.400 2.635 ;
        RECT 0.570 1.665 0.820 2.465 ;
        RECT 0.990 1.835 1.770 2.635 ;
        RECT 0.570 1.495 1.340 1.665 ;
        RECT 1.170 1.325 1.340 1.495 ;
        RECT 2.820 1.455 3.070 2.635 ;
        RECT 1.170 0.995 1.470 1.325 ;
        RECT 1.170 0.825 1.340 0.995 ;
        RECT 0.090 0.085 0.425 0.815 ;
        RECT 1.000 0.280 1.340 0.825 ;
        RECT 1.980 0.725 3.110 0.905 ;
        RECT 1.980 0.425 2.270 0.725 ;
        RECT 2.440 0.085 2.610 0.555 ;
        RECT 2.780 0.275 3.110 0.725 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__o2bb2ai_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o2bb2ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.445 1.945 1.615 ;
        RECT 0.090 1.075 0.625 1.445 ;
        RECT 1.615 1.075 1.945 1.445 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.795 1.075 1.400 1.275 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.410 1.445 5.435 1.615 ;
        RECT 3.410 1.075 3.740 1.445 ;
        RECT 4.730 1.075 5.435 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.960 1.075 4.500 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.300 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.715500 ;
    PORT
      LAYER li1 ;
        RECT 2.745 1.955 3.035 2.465 ;
        RECT 4.080 1.955 4.330 2.125 ;
        RECT 2.745 1.785 4.330 1.955 ;
        RECT 2.745 1.075 3.215 1.785 ;
        RECT 2.745 0.645 3.075 1.075 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.150 1.795 0.400 2.635 ;
        RECT 0.575 1.965 0.825 2.465 ;
        RECT 0.995 2.135 1.245 2.635 ;
        RECT 1.835 2.135 2.575 2.635 ;
        RECT 3.205 2.125 3.490 2.635 ;
        RECT 3.660 2.295 4.750 2.465 ;
        RECT 3.660 2.125 3.910 2.295 ;
        RECT 1.415 1.965 1.665 2.125 ;
        RECT 0.575 1.785 2.285 1.965 ;
        RECT 4.500 1.785 4.750 2.295 ;
        RECT 4.965 1.795 5.170 2.635 ;
        RECT 2.115 1.325 2.285 1.785 ;
        RECT 2.115 0.995 2.575 1.325 ;
        RECT 2.115 0.905 2.285 0.995 ;
        RECT 0.195 0.085 0.365 0.895 ;
        RECT 0.535 0.475 0.785 0.895 ;
        RECT 0.955 0.725 2.285 0.905 ;
        RECT 3.245 0.735 5.210 0.905 ;
        RECT 0.955 0.645 1.285 0.725 ;
        RECT 0.535 0.305 1.705 0.475 ;
        RECT 1.875 0.085 2.045 0.555 ;
        RECT 2.325 0.475 2.575 0.555 ;
        RECT 3.245 0.475 3.530 0.735 ;
        RECT 4.040 0.725 5.210 0.735 ;
        RECT 2.325 0.255 3.530 0.475 ;
        RECT 3.700 0.085 3.870 0.555 ;
        RECT 4.040 0.255 4.370 0.725 ;
        RECT 4.540 0.085 4.710 0.555 ;
        RECT 4.880 0.255 5.210 0.725 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__o2bb2ai_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o2bb2ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2bb2ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 2.095 1.075 3.505 1.285 ;
    END
  END A1_N
  PIN A2_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.075 1.825 1.285 ;
    END
  END A2_N
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 8.045 1.075 10.005 1.285 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.465 1.075 7.875 1.285 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.945 1.015 ;
        RECT 0.135 -0.085 0.305 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.431000 ;
    PORT
      LAYER li1 ;
        RECT 4.425 1.625 4.675 2.465 ;
        RECT 5.265 1.625 5.515 2.465 ;
        RECT 6.625 1.625 6.875 2.125 ;
        RECT 7.465 1.625 7.715 2.125 ;
        RECT 4.425 1.455 7.715 1.625 ;
        RECT 5.875 0.905 6.155 1.455 ;
        RECT 4.415 0.645 6.155 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.155 1.795 0.405 2.635 ;
        RECT 0.575 1.625 0.825 2.465 ;
        RECT 0.995 1.795 1.245 2.635 ;
        RECT 1.415 1.625 1.665 2.465 ;
        RECT 1.835 1.795 2.085 2.635 ;
        RECT 2.255 1.625 2.505 2.465 ;
        RECT 2.675 1.795 2.925 2.635 ;
        RECT 3.095 1.625 3.345 2.465 ;
        RECT 3.515 1.795 4.255 2.635 ;
        RECT 4.845 1.795 5.095 2.635 ;
        RECT 5.685 1.795 5.935 2.635 ;
        RECT 6.175 2.295 8.135 2.465 ;
        RECT 6.175 1.795 6.455 2.295 ;
        RECT 7.045 1.795 7.295 2.295 ;
        RECT 7.885 1.625 8.135 2.295 ;
        RECT 8.305 1.795 8.555 2.635 ;
        RECT 8.725 1.625 8.975 2.465 ;
        RECT 9.145 1.795 9.395 2.635 ;
        RECT 9.565 1.625 9.875 2.465 ;
        RECT 0.085 1.455 3.915 1.625 ;
        RECT 7.885 1.455 9.875 1.625 ;
        RECT 0.085 0.905 0.255 1.455 ;
        RECT 3.745 1.285 3.915 1.455 ;
        RECT 3.745 1.075 5.705 1.285 ;
        RECT 0.085 0.645 1.705 0.905 ;
        RECT 1.875 0.725 3.805 0.905 ;
        RECT 1.875 0.475 2.125 0.725 ;
        RECT 0.100 0.255 2.125 0.475 ;
        RECT 2.295 0.085 2.465 0.555 ;
        RECT 2.635 0.255 2.965 0.725 ;
        RECT 3.135 0.085 3.305 0.555 ;
        RECT 3.475 0.255 3.805 0.725 ;
        RECT 4.060 0.475 4.245 0.835 ;
        RECT 6.325 0.735 9.855 0.905 ;
        RECT 6.325 0.475 6.495 0.735 ;
        RECT 7.005 0.725 9.855 0.735 ;
        RECT 4.060 0.255 6.495 0.475 ;
        RECT 6.665 0.085 6.835 0.555 ;
        RECT 7.005 0.255 7.335 0.725 ;
        RECT 7.505 0.085 7.675 0.555 ;
        RECT 7.845 0.255 8.175 0.725 ;
        RECT 8.345 0.085 8.515 0.555 ;
        RECT 8.685 0.255 9.015 0.725 ;
        RECT 9.185 0.085 9.355 0.555 ;
        RECT 9.525 0.255 9.855 0.725 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
  END
END sky130_fd_sc_hd__o2bb2ai_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o21a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.275 2.675 1.615 ;
        RECT 2.345 1.075 2.675 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.940 1.275 2.155 2.390 ;
        RECT 1.705 1.095 2.155 1.275 ;
        RECT 1.705 1.075 2.035 1.095 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.075 1.535 1.305 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.755 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.449000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.030 0.365 2.465 ;
        RECT 0.085 0.255 0.425 1.030 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.535 1.860 1.245 2.635 ;
        RECT 1.415 1.690 1.745 2.465 ;
        RECT 2.335 1.915 2.665 2.635 ;
        RECT 0.595 1.475 1.745 1.690 ;
        RECT 0.595 0.905 0.880 1.475 ;
        RECT 0.595 0.715 1.305 0.905 ;
        RECT 1.005 0.575 1.305 0.715 ;
        RECT 1.495 0.715 2.675 0.905 ;
        RECT 1.495 0.635 1.825 0.715 ;
        RECT 1.005 0.565 1.320 0.575 ;
        RECT 1.005 0.555 1.330 0.565 ;
        RECT 1.005 0.550 1.340 0.555 ;
        RECT 0.595 0.085 0.765 0.545 ;
        RECT 1.005 0.540 1.345 0.550 ;
        RECT 1.005 0.535 1.350 0.540 ;
        RECT 1.005 0.525 1.355 0.535 ;
        RECT 1.005 0.520 1.360 0.525 ;
        RECT 1.005 0.255 1.365 0.520 ;
        RECT 1.995 0.085 2.165 0.545 ;
        RECT 2.335 0.255 2.675 0.715 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__o21a_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o21a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.865 0.995 3.125 1.450 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.400 2.610 1.985 ;
        RECT 2.025 1.025 2.610 1.400 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.445 1.010 1.855 1.615 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.215 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.453750 ;
    PORT
      LAYER li1 ;
        RECT 0.530 0.255 0.775 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.090 1.635 0.345 2.635 ;
        RECT 0.945 2.185 1.795 2.635 ;
        RECT 1.965 2.005 2.225 2.465 ;
        RECT 1.105 1.785 2.225 2.005 ;
        RECT 1.105 1.330 1.275 1.785 ;
        RECT 2.795 1.650 3.120 2.635 ;
        RECT 0.105 0.085 0.345 0.885 ;
        RECT 0.945 0.840 1.275 1.330 ;
        RECT 0.945 0.635 1.795 0.840 ;
        RECT 0.945 0.085 1.275 0.465 ;
        RECT 1.465 0.255 1.795 0.635 ;
        RECT 1.965 0.635 3.120 0.825 ;
        RECT 1.965 0.465 2.175 0.635 ;
        RECT 2.845 0.495 3.120 0.635 ;
        RECT 2.345 0.085 2.675 0.465 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__o21a_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o21a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.480 1.495 5.400 1.705 ;
        RECT 3.480 0.990 3.785 1.495 ;
        RECT 5.030 0.995 5.400 1.495 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.140 0.995 4.690 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.485 1.075 3.155 1.615 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.495 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.924000 ;
    PORT
      LAYER li1 ;
        RECT 0.915 1.700 1.105 2.465 ;
        RECT 1.775 1.700 1.955 2.465 ;
        RECT 0.090 1.530 1.955 1.700 ;
        RECT 0.090 0.805 0.320 1.530 ;
        RECT 0.090 0.635 1.715 0.805 ;
        RECT 0.595 0.615 1.715 0.635 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.415 1.870 0.745 2.635 ;
        RECT 1.275 1.870 1.605 2.635 ;
        RECT 2.135 2.255 2.485 2.635 ;
        RECT 2.655 2.105 2.845 2.465 ;
        RECT 3.015 2.275 3.685 2.635 ;
        RECT 4.215 2.105 4.545 2.445 ;
        RECT 2.655 2.085 4.545 2.105 ;
        RECT 2.125 1.875 4.545 2.085 ;
        RECT 5.075 1.935 5.435 2.635 ;
        RECT 2.125 1.830 2.845 1.875 ;
        RECT 2.125 1.335 2.315 1.830 ;
        RECT 0.490 0.995 2.315 1.335 ;
        RECT 2.115 0.870 2.315 0.995 ;
        RECT 2.115 0.655 3.095 0.870 ;
        RECT 3.275 0.615 5.405 0.785 ;
        RECT 3.275 0.485 3.605 0.615 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 0.955 0.085 1.285 0.445 ;
        RECT 1.815 0.085 2.145 0.465 ;
        RECT 2.335 0.255 3.605 0.485 ;
        RECT 3.775 0.085 4.115 0.445 ;
        RECT 4.645 0.085 4.975 0.445 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__o21a_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o21ai_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.415 1.615 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.340 0.775 1.645 ;
        RECT 0.605 1.100 1.005 1.340 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.355 1.730 1.685 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.105 1.830 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.290500 ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.680 1.300 2.465 ;
        RECT 0.965 1.510 1.345 1.680 ;
        RECT 1.175 1.125 1.345 1.510 ;
        RECT 1.175 0.955 1.740 1.125 ;
        RECT 1.455 0.280 1.740 0.955 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.145 1.825 0.475 2.635 ;
        RECT 1.470 1.855 1.725 2.635 ;
        RECT 0.120 0.615 1.285 0.785 ;
        RECT 0.120 0.280 0.380 0.615 ;
        RECT 0.550 0.085 0.880 0.445 ;
        RECT 1.050 0.280 1.285 0.615 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__o21ai_0

#--------EOF---------

MACRO sky130_fd_sc_hd__o21ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.150 0.995 0.410 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.590 1.325 0.785 2.375 ;
        RECT 0.590 0.995 0.975 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.202500 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.295 1.750 1.655 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 1.840 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 1.835 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.030 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 1.840 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.517000 ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.785 1.295 2.465 ;
        RECT 0.965 1.505 1.315 1.785 ;
        RECT 1.145 1.125 1.315 1.505 ;
        RECT 1.145 0.955 1.665 1.125 ;
        RECT 1.495 0.390 1.665 0.955 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 1.840 2.805 ;
        RECT 0.090 1.495 0.410 2.635 ;
        RECT 1.495 1.835 1.750 2.635 ;
        RECT 0.090 0.615 1.305 0.785 ;
        RECT 0.090 0.265 0.380 0.615 ;
        RECT 0.575 0.085 0.905 0.445 ;
        RECT 1.075 0.310 1.305 0.615 ;
        RECT 0.000 -0.085 1.840 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
  END
END sky130_fd_sc_hd__o21ai_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o21ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.120 1.445 2.095 1.615 ;
        RECT 0.120 1.055 0.450 1.445 ;
        RECT 1.600 1.075 2.095 1.445 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.620 1.075 1.420 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.815 0.765 3.130 1.400 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.105 3.215 1.015 ;
        RECT 0.140 -0.085 0.310 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.742000 ;
    PORT
      LAYER li1 ;
        RECT 0.995 1.965 1.295 2.125 ;
        RECT 2.410 1.965 2.645 2.465 ;
        RECT 0.995 1.785 2.645 1.965 ;
        RECT 2.435 0.595 2.645 1.785 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.105 1.785 0.435 2.635 ;
        RECT 0.605 2.295 1.715 2.465 ;
        RECT 0.605 1.785 0.825 2.295 ;
        RECT 1.525 2.135 1.715 2.295 ;
        RECT 1.910 2.175 2.240 2.635 ;
        RECT 2.815 1.570 3.125 2.635 ;
        RECT 0.105 0.715 2.265 0.885 ;
        RECT 0.105 0.255 0.435 0.715 ;
        RECT 0.615 0.085 0.785 0.545 ;
        RECT 0.965 0.255 1.295 0.715 ;
        RECT 1.525 0.085 1.695 0.545 ;
        RECT 1.935 0.425 2.265 0.715 ;
        RECT 2.815 0.425 3.125 0.595 ;
        RECT 1.935 0.255 3.125 0.425 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__o21ai_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o21ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.575 1.515 3.695 1.685 ;
        RECT 0.575 1.320 1.475 1.515 ;
        RECT 0.125 1.015 1.475 1.320 ;
        RECT 3.445 0.990 3.695 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.985 1.070 3.275 1.345 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.905 1.015 5.255 1.275 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.105 5.760 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.484000 ;
    PORT
      LAYER li1 ;
        RECT 4.080 2.085 4.290 2.465 ;
        RECT 4.960 2.085 5.150 2.465 ;
        RECT 4.080 2.025 5.150 2.085 ;
        RECT 1.840 1.855 5.150 2.025 ;
        RECT 3.935 1.700 5.150 1.855 ;
        RECT 3.935 1.445 5.835 1.700 ;
        RECT 5.425 0.845 5.835 1.445 ;
        RECT 4.030 0.615 5.835 0.845 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.120 1.820 0.405 2.635 ;
        RECT 0.575 2.085 0.810 2.465 ;
        RECT 0.980 2.255 1.310 2.635 ;
        RECT 1.480 2.275 3.460 2.465 ;
        RECT 1.480 2.085 1.670 2.275 ;
        RECT 3.630 2.195 3.910 2.635 ;
        RECT 4.460 2.255 4.790 2.635 ;
        RECT 0.575 1.915 1.670 2.085 ;
        RECT 5.320 1.880 5.650 2.635 ;
        RECT 0.120 0.615 3.860 0.820 ;
        RECT 3.630 0.445 3.860 0.615 ;
        RECT 0.550 0.085 0.880 0.445 ;
        RECT 1.410 0.085 1.740 0.445 ;
        RECT 2.270 0.085 2.600 0.445 ;
        RECT 3.130 0.085 3.460 0.445 ;
        RECT 3.630 0.255 5.650 0.445 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
END sky130_fd_sc_hd__o21ai_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o21ba_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ba_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.950 1.075 3.595 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.210 1.075 2.780 1.285 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.030 0.995 1.360 1.325 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.085 0.105 3.535 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.480 0.425 2.465 ;
        RECT 0.085 0.825 0.340 1.480 ;
        RECT 0.085 0.450 0.445 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.595 2.205 1.005 2.635 ;
        RECT 1.750 2.215 2.080 2.635 ;
        RECT 2.250 2.035 2.575 2.465 ;
        RECT 0.595 1.865 2.575 2.035 ;
        RECT 0.595 1.325 0.860 1.865 ;
        RECT 1.075 1.525 1.700 1.695 ;
        RECT 0.510 0.995 0.860 1.325 ;
        RECT 1.530 0.825 1.700 1.525 ;
        RECT 0.710 0.085 0.880 0.825 ;
        RECT 1.160 0.655 1.700 0.825 ;
        RECT 1.870 1.455 2.575 1.865 ;
        RECT 3.050 1.535 3.380 2.635 ;
        RECT 1.160 0.450 1.330 0.655 ;
        RECT 1.870 0.255 2.040 1.455 ;
        RECT 2.270 0.735 3.440 0.905 ;
        RECT 2.270 0.255 2.600 0.735 ;
        RECT 2.770 0.085 2.940 0.555 ;
        RECT 3.110 0.270 3.440 0.735 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__o21ba_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o21ba_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ba_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.100 1.075 3.595 1.625 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.075 2.930 1.285 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.325 0.775 1.695 ;
        RECT 0.425 0.995 0.775 1.325 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 3.675 1.015 ;
        RECT 0.145 0.105 3.675 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.945 1.495 1.350 1.695 ;
        RECT 0.945 0.595 1.115 1.495 ;
        RECT 0.945 0.255 1.240 0.595 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.520 2.205 0.910 2.635 ;
        RECT 1.415 2.205 2.230 2.635 ;
        RECT 2.400 2.035 2.725 2.465 ;
        RECT 0.085 1.865 1.935 2.035 ;
        RECT 0.085 1.495 0.395 1.865 ;
        RECT 0.085 0.825 0.255 1.495 ;
        RECT 1.285 1.060 1.455 1.325 ;
        RECT 1.285 0.890 1.595 1.060 ;
        RECT 1.765 0.995 1.935 1.865 ;
        RECT 2.105 1.455 2.725 2.035 ;
        RECT 3.200 1.875 3.530 2.635 ;
        RECT 1.425 0.825 1.595 0.890 ;
        RECT 2.105 0.825 2.275 1.455 ;
        RECT 0.085 0.430 0.345 0.825 ;
        RECT 0.595 0.085 0.775 0.825 ;
        RECT 1.425 0.655 2.275 0.825 ;
        RECT 1.410 0.085 1.770 0.485 ;
        RECT 1.940 0.255 2.275 0.655 ;
        RECT 2.445 0.735 3.590 0.905 ;
        RECT 2.445 0.365 2.745 0.735 ;
        RECT 2.915 0.085 3.085 0.555 ;
        RECT 3.255 0.270 3.590 0.735 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__o21ba_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o21ba_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21ba_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.990 1.075 5.895 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.780 1.075 4.820 1.275 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.285 0.885 1.705 ;
        RECT 0.425 1.075 0.885 1.285 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.080 0.105 5.795 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 1.055 1.445 2.225 1.705 ;
        RECT 1.055 0.905 1.455 1.445 ;
        RECT 1.055 0.725 2.225 0.905 ;
        RECT 1.055 0.255 1.385 0.725 ;
        RECT 1.895 0.255 2.225 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.085 2.045 0.435 2.465 ;
        RECT 0.635 2.215 0.965 2.635 ;
        RECT 1.475 2.215 1.805 2.635 ;
        RECT 2.315 2.215 2.645 2.635 ;
        RECT 0.085 1.875 2.565 2.045 ;
        RECT 0.085 1.455 0.435 1.875 ;
        RECT 2.395 1.615 2.565 1.875 ;
        RECT 2.815 1.965 2.985 2.465 ;
        RECT 3.200 2.135 3.450 2.635 ;
        RECT 3.685 2.295 4.765 2.465 ;
        RECT 3.685 2.135 3.925 2.295 ;
        RECT 4.135 1.965 4.380 2.125 ;
        RECT 2.815 1.795 4.380 1.965 ;
        RECT 0.085 0.855 0.255 1.455 ;
        RECT 2.395 1.445 2.905 1.615 ;
        RECT 1.625 1.075 2.565 1.275 ;
        RECT 2.735 1.245 2.905 1.445 ;
        RECT 2.735 1.075 3.135 1.245 ;
        RECT 0.085 0.265 0.545 0.855 ;
        RECT 0.715 0.085 0.885 0.905 ;
        RECT 2.395 0.895 2.565 1.075 ;
        RECT 3.395 0.895 3.585 1.795 ;
        RECT 4.135 1.445 4.380 1.795 ;
        RECT 4.595 1.665 4.765 2.295 ;
        RECT 4.935 1.835 5.265 2.635 ;
        RECT 5.435 1.665 5.710 2.465 ;
        RECT 4.595 1.455 5.710 1.665 ;
        RECT 2.395 0.725 3.585 0.895 ;
        RECT 3.235 0.645 3.585 0.725 ;
        RECT 3.755 0.725 5.710 0.905 ;
        RECT 1.555 0.085 1.725 0.555 ;
        RECT 2.395 0.085 2.565 0.555 ;
        RECT 3.755 0.475 4.005 0.725 ;
        RECT 2.805 0.255 4.005 0.475 ;
        RECT 4.175 0.085 4.345 0.555 ;
        RECT 4.515 0.255 4.845 0.725 ;
        RECT 5.015 0.085 5.185 0.555 ;
        RECT 5.355 0.265 5.710 0.725 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
END sky130_fd_sc_hd__o21ba_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o21bai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21bai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.195 1.075 2.675 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.075 2.025 1.285 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.345 0.355 2.445 ;
        RECT 0.085 0.995 0.535 1.345 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 2.755 1.015 ;
        RECT 0.145 0.105 2.755 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.474000 ;
    PORT
      LAYER li1 ;
        RECT 1.470 1.625 1.795 2.465 ;
        RECT 1.185 1.455 1.795 1.625 ;
        RECT 1.185 0.825 1.355 1.455 ;
        RECT 1.115 0.645 1.355 0.825 ;
        RECT 1.115 0.255 1.285 0.645 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.525 1.705 0.800 2.210 ;
        RECT 0.970 1.875 1.300 2.635 ;
        RECT 0.525 1.535 1.015 1.705 ;
        RECT 2.270 1.535 2.645 2.635 ;
        RECT 0.720 0.995 1.015 1.535 ;
        RECT 0.720 0.825 0.890 0.995 ;
        RECT 0.085 0.085 0.360 0.825 ;
        RECT 0.580 0.655 0.890 0.825 ;
        RECT 1.570 0.735 2.665 0.905 ;
        RECT 0.580 0.495 0.770 0.655 ;
        RECT 1.570 0.485 1.740 0.735 ;
        RECT 1.490 0.255 1.820 0.485 ;
        RECT 1.995 0.085 2.165 0.555 ;
        RECT 2.335 0.270 2.665 0.735 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__o21bai_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o21bai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21bai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.260 1.075 4.055 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.950 1.075 3.090 1.275 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.525 1.325 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.335 4.065 1.015 ;
        RECT 0.145 0.105 4.065 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.715500 ;
    PORT
      LAYER li1 ;
        RECT 1.085 1.615 1.255 2.465 ;
        RECT 2.405 1.615 2.650 2.125 ;
        RECT 1.085 1.445 2.650 1.615 ;
        RECT 1.525 0.905 1.780 1.445 ;
        RECT 1.525 0.645 1.855 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.180 1.665 0.350 1.915 ;
        RECT 0.585 1.875 0.915 2.635 ;
        RECT 1.470 1.795 1.720 2.635 ;
        RECT 1.955 2.295 3.035 2.465 ;
        RECT 1.955 1.795 2.235 2.295 ;
        RECT 2.865 1.665 3.035 2.295 ;
        RECT 3.205 1.835 3.535 2.635 ;
        RECT 3.705 1.665 3.980 2.465 ;
        RECT 0.180 1.495 0.865 1.665 ;
        RECT 0.695 1.245 0.865 1.495 ;
        RECT 2.865 1.455 3.980 1.665 ;
        RECT 0.695 1.075 1.335 1.245 ;
        RECT 0.695 0.825 0.865 1.075 ;
        RECT 0.180 0.085 0.350 0.825 ;
        RECT 0.600 0.445 0.865 0.825 ;
        RECT 1.075 0.475 1.355 0.905 ;
        RECT 2.025 0.725 3.980 0.905 ;
        RECT 2.025 0.475 2.275 0.725 ;
        RECT 1.075 0.255 2.275 0.475 ;
        RECT 2.445 0.085 2.615 0.555 ;
        RECT 2.785 0.255 3.115 0.725 ;
        RECT 3.285 0.085 3.455 0.555 ;
        RECT 3.625 0.265 3.980 0.725 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__o21bai_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o21bai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o21bai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.585 1.285 6.810 2.455 ;
        RECT 4.645 1.075 6.810 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.065 1.075 4.475 1.275 ;
    END
  END A2
  PIN B1_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.555 1.285 ;
    END
  END B1_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.035 0.105 6.545 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.431000 ;
    PORT
      LAYER li1 ;
        RECT 1.065 1.625 1.275 2.465 ;
        RECT 1.865 1.625 2.115 2.465 ;
        RECT 3.225 1.625 3.475 2.125 ;
        RECT 4.065 1.625 4.315 2.125 ;
        RECT 1.065 1.455 4.315 1.625 ;
        RECT 2.445 1.445 4.315 1.455 ;
        RECT 2.445 1.075 2.895 1.445 ;
        RECT 2.445 0.815 2.675 1.075 ;
        RECT 1.420 0.645 2.675 0.815 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.145 1.625 0.475 2.435 ;
        RECT 0.645 1.795 0.855 2.635 ;
        RECT 1.445 1.795 1.695 2.635 ;
        RECT 2.285 1.795 2.535 2.635 ;
        RECT 2.775 2.295 4.735 2.465 ;
        RECT 2.775 1.795 3.055 2.295 ;
        RECT 3.645 1.795 3.895 2.295 ;
        RECT 4.485 1.625 4.735 2.295 ;
        RECT 4.905 1.795 5.155 2.635 ;
        RECT 5.325 1.625 5.575 2.465 ;
        RECT 5.745 1.795 5.995 2.635 ;
        RECT 6.165 1.625 6.415 2.465 ;
        RECT 0.145 1.455 0.895 1.625 ;
        RECT 4.485 1.455 6.415 1.625 ;
        RECT 0.725 1.285 0.895 1.455 ;
        RECT 0.725 1.075 2.275 1.285 ;
        RECT 0.725 0.895 0.895 1.075 ;
        RECT 0.225 0.085 0.395 0.895 ;
        RECT 0.565 0.290 0.895 0.895 ;
        RECT 2.845 0.725 6.455 0.905 ;
        RECT 2.845 0.475 3.095 0.725 ;
        RECT 1.080 0.305 3.095 0.475 ;
        RECT 3.265 0.085 3.435 0.555 ;
        RECT 3.605 0.255 3.935 0.725 ;
        RECT 4.105 0.085 4.275 0.555 ;
        RECT 4.445 0.255 4.775 0.725 ;
        RECT 4.945 0.085 5.115 0.555 ;
        RECT 5.285 0.255 5.615 0.725 ;
        RECT 5.785 0.085 5.955 0.555 ;
        RECT 6.125 0.255 6.455 0.725 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
  END
END sky130_fd_sc_hd__o21bai_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o22a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.670 1.075 3.135 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.615 2.645 2.405 ;
        RECT 2.315 1.445 2.645 1.615 ;
        RECT 2.315 1.325 2.495 1.445 ;
        RECT 2.165 1.075 2.495 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.980 1.075 1.335 1.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.530 1.075 1.995 1.325 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.215 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.449000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.365 0.365 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.555 1.875 1.340 2.635 ;
        RECT 1.735 1.805 2.120 2.465 ;
        RECT 1.735 1.705 2.145 1.805 ;
        RECT 0.535 1.495 2.145 1.705 ;
        RECT 0.535 0.895 0.810 1.495 ;
        RECT 2.815 1.455 3.135 2.635 ;
        RECT 0.535 0.715 1.785 0.895 ;
        RECT 1.420 0.645 1.785 0.715 ;
        RECT 1.955 0.695 3.135 0.865 ;
        RECT 0.595 0.085 0.765 0.545 ;
        RECT 1.955 0.475 2.285 0.695 ;
        RECT 1.035 0.295 2.285 0.475 ;
        RECT 2.455 0.085 2.625 0.525 ;
        RECT 2.795 0.280 3.135 0.695 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__o22a_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o22a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.270 1.275 3.590 1.615 ;
        RECT 3.095 1.075 3.590 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.900 1.615 3.100 2.405 ;
        RECT 2.745 1.445 3.100 1.615 ;
        RECT 2.745 1.325 2.925 1.445 ;
        RECT 2.595 1.075 2.925 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.435 1.075 1.790 1.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.960 1.075 2.425 1.325 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.105 3.675 1.015 ;
        RECT 0.130 -0.085 0.300 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.590 0.365 0.805 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.115 1.445 0.365 2.635 ;
        RECT 0.995 1.875 1.795 2.635 ;
        RECT 2.190 1.705 2.575 2.465 ;
        RECT 3.270 1.795 3.590 2.635 ;
        RECT 0.975 1.495 2.575 1.705 ;
        RECT 0.975 0.895 1.255 1.495 ;
        RECT 0.185 0.085 0.355 0.885 ;
        RECT 0.975 0.715 2.215 0.895 ;
        RECT 2.560 0.825 3.590 0.865 ;
        RECT 1.850 0.645 2.215 0.715 ;
        RECT 2.390 0.695 3.590 0.825 ;
        RECT 1.025 0.085 1.205 0.545 ;
        RECT 2.390 0.475 2.730 0.695 ;
        RECT 1.465 0.295 2.730 0.475 ;
        RECT 2.915 0.085 3.085 0.525 ;
        RECT 3.255 0.280 3.590 0.695 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__o22a_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o22a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.350 1.445 5.735 1.615 ;
        RECT 4.350 1.075 4.680 1.445 ;
        RECT 5.565 1.275 5.735 1.445 ;
        RECT 5.565 1.075 6.355 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.900 1.075 5.395 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.420 1.445 4.180 1.615 ;
        RECT 2.420 1.075 2.955 1.445 ;
        RECT 3.850 1.075 4.180 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.125 1.075 3.680 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.070 0.105 6.240 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.640 1.615 0.890 2.465 ;
        RECT 1.480 1.615 1.730 2.465 ;
        RECT 0.085 1.445 1.730 1.615 ;
        RECT 0.085 0.905 0.370 1.445 ;
        RECT 0.085 0.725 1.770 0.905 ;
        RECT 0.600 0.265 0.930 0.725 ;
        RECT 1.440 0.255 1.770 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.220 1.825 0.470 2.635 ;
        RECT 1.060 1.795 1.310 2.635 ;
        RECT 1.900 2.125 2.670 2.635 ;
        RECT 2.840 2.295 3.930 2.465 ;
        RECT 2.840 2.125 3.090 2.295 ;
        RECT 3.680 2.125 3.930 2.295 ;
        RECT 4.100 2.125 4.430 2.635 ;
        RECT 4.600 2.295 5.690 2.465 ;
        RECT 4.600 2.125 4.850 2.295 ;
        RECT 3.260 1.955 3.510 2.125 ;
        RECT 5.020 1.955 5.270 2.125 ;
        RECT 1.900 1.785 5.270 1.955 ;
        RECT 5.440 1.785 5.690 2.295 ;
        RECT 1.900 1.275 2.230 1.785 ;
        RECT 5.905 1.455 6.110 2.635 ;
        RECT 0.540 1.075 2.230 1.275 ;
        RECT 1.940 0.905 2.230 1.075 ;
        RECT 1.940 0.735 3.970 0.905 ;
        RECT 2.415 0.645 3.970 0.735 ;
        RECT 4.140 0.735 6.150 0.905 ;
        RECT 0.260 0.085 0.430 0.555 ;
        RECT 1.100 0.085 1.270 0.555 ;
        RECT 1.940 0.085 2.110 0.555 ;
        RECT 4.140 0.475 4.470 0.735 ;
        RECT 4.980 0.725 6.150 0.735 ;
        RECT 2.380 0.255 4.470 0.475 ;
        RECT 4.640 0.085 4.810 0.555 ;
        RECT 4.980 0.255 5.310 0.725 ;
        RECT 5.480 0.085 5.650 0.555 ;
        RECT 5.820 0.255 6.150 0.725 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
END sky130_fd_sc_hd__o22a_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o22ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.755 1.075 2.215 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.615 1.725 2.405 ;
        RECT 1.405 1.445 1.725 1.615 ;
        RECT 1.405 1.245 1.585 1.445 ;
        RECT 1.220 1.075 1.585 1.245 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.665 0.325 1.990 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.835 1.415 1.235 1.665 ;
        RECT 0.835 0.995 1.005 1.415 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.295 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.650250 ;
    PORT
      LAYER li1 ;
        RECT 0.835 2.045 1.335 2.465 ;
        RECT 0.495 1.835 1.335 2.045 ;
        RECT 0.495 0.825 0.665 1.835 ;
        RECT 0.495 0.645 0.845 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.135 2.175 0.345 2.635 ;
        RECT 1.895 1.455 2.215 2.635 ;
        RECT 1.185 0.825 2.215 0.865 ;
        RECT 1.015 0.695 2.215 0.825 ;
        RECT 1.015 0.475 1.345 0.695 ;
        RECT 0.085 0.295 1.345 0.475 ;
        RECT 1.535 0.085 1.705 0.525 ;
        RECT 1.875 0.280 2.215 0.695 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__o22ai_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o22ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.075 4.165 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.555 1.075 3.225 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.200 1.075 0.985 1.285 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.155 1.075 1.925 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.455 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 1.415 1.625 1.665 2.125 ;
        RECT 2.815 1.625 3.065 2.125 ;
        RECT 1.415 1.445 3.065 1.625 ;
        RECT 2.095 0.905 2.340 1.445 ;
        RECT 0.535 0.725 2.340 0.905 ;
        RECT 0.535 0.645 0.865 0.725 ;
        RECT 1.375 0.645 1.705 0.725 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.150 1.625 0.405 2.465 ;
        RECT 0.575 1.795 0.825 2.635 ;
        RECT 0.995 2.295 2.085 2.465 ;
        RECT 0.995 1.625 1.245 2.295 ;
        RECT 1.835 1.795 2.085 2.295 ;
        RECT 2.395 2.295 3.485 2.465 ;
        RECT 2.395 1.795 2.645 2.295 ;
        RECT 0.150 1.455 1.245 1.625 ;
        RECT 3.235 1.625 3.485 2.295 ;
        RECT 3.655 1.795 3.905 2.635 ;
        RECT 4.075 1.625 4.330 2.465 ;
        RECT 3.235 1.455 4.330 1.625 ;
        RECT 0.090 0.475 0.365 0.905 ;
        RECT 2.510 0.725 4.365 0.905 ;
        RECT 2.510 0.475 2.680 0.725 ;
        RECT 0.090 0.305 2.680 0.475 ;
        RECT 2.855 0.085 3.025 0.555 ;
        RECT 3.195 0.255 3.525 0.725 ;
        RECT 3.695 0.085 3.865 0.555 ;
        RECT 4.035 0.255 4.365 0.725 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__o22ai_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o22ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o22ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.150 1.445 3.575 1.615 ;
        RECT 1.150 1.275 1.415 1.445 ;
        RECT 0.085 1.075 1.415 1.275 ;
        RECT 3.275 1.245 3.575 1.445 ;
        RECT 3.275 1.075 3.605 1.245 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.685 1.075 3.095 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 4.295 1.445 6.935 1.615 ;
        RECT 4.295 0.995 4.940 1.445 ;
        RECT 6.715 0.995 6.935 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 5.110 1.075 6.460 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.035 0.105 7.315 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 1.845 1.955 2.095 2.125 ;
        RECT 2.685 1.955 2.935 2.125 ;
        RECT 5.255 1.955 5.505 2.125 ;
        RECT 6.095 1.955 6.345 2.125 ;
        RECT 1.845 1.785 3.915 1.955 ;
        RECT 5.255 1.785 7.275 1.955 ;
        RECT 3.745 1.615 3.915 1.785 ;
        RECT 3.745 1.445 4.125 1.615 ;
        RECT 3.955 0.820 4.125 1.445 ;
        RECT 7.105 0.820 7.275 1.785 ;
        RECT 3.955 0.645 7.275 0.820 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.165 1.445 0.415 2.635 ;
        RECT 0.585 1.955 0.835 2.465 ;
        RECT 1.005 2.125 1.255 2.635 ;
        RECT 1.425 2.295 3.395 2.465 ;
        RECT 1.425 1.955 1.675 2.295 ;
        RECT 2.265 2.125 2.515 2.295 ;
        RECT 3.105 2.125 3.395 2.295 ;
        RECT 3.565 2.125 3.785 2.635 ;
        RECT 3.955 2.125 4.255 2.465 ;
        RECT 4.425 2.125 4.665 2.635 ;
        RECT 4.835 2.295 6.765 2.465 ;
        RECT 0.585 1.785 1.675 1.955 ;
        RECT 4.085 1.955 4.255 2.125 ;
        RECT 4.835 1.955 5.085 2.295 ;
        RECT 5.675 2.125 5.925 2.295 ;
        RECT 6.515 2.135 6.765 2.295 ;
        RECT 6.935 2.125 7.215 2.635 ;
        RECT 4.085 1.785 5.085 1.955 ;
        RECT 0.585 1.445 0.835 1.785 ;
        RECT 0.125 0.735 3.785 0.905 ;
        RECT 0.125 0.725 1.295 0.735 ;
        RECT 0.125 0.255 0.455 0.725 ;
        RECT 0.625 0.085 0.795 0.555 ;
        RECT 0.965 0.255 1.295 0.725 ;
        RECT 1.805 0.725 2.975 0.735 ;
        RECT 1.465 0.085 1.635 0.555 ;
        RECT 1.805 0.255 2.135 0.725 ;
        RECT 2.305 0.085 2.475 0.555 ;
        RECT 2.645 0.255 2.975 0.725 ;
        RECT 3.145 0.085 3.315 0.555 ;
        RECT 3.485 0.475 3.785 0.735 ;
        RECT 3.485 0.255 7.245 0.475 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
END sky130_fd_sc_hd__o22ai_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o31a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.905 0.995 1.295 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.325 1.725 2.125 ;
        RECT 1.480 0.995 1.725 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.925 0.995 2.175 2.125 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.390 0.995 2.795 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.085 0.105 3.085 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.594000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.835 0.525 2.465 ;
        RECT 0.085 0.825 0.395 1.835 ;
        RECT 0.085 0.265 0.525 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.700 1.785 1.015 2.635 ;
        RECT 1.185 2.295 2.615 2.465 ;
        RECT 1.185 1.615 1.355 2.295 ;
        RECT 0.565 1.445 1.355 1.615 ;
        RECT 2.365 1.665 2.615 2.295 ;
        RECT 2.795 1.835 3.125 2.635 ;
        RECT 2.365 1.495 3.135 1.665 ;
        RECT 0.565 0.995 0.735 1.445 ;
        RECT 2.965 0.825 3.135 1.495 ;
        RECT 0.695 0.085 1.145 0.825 ;
        RECT 1.315 0.655 2.475 0.825 ;
        RECT 1.315 0.255 1.485 0.655 ;
        RECT 1.655 0.085 2.075 0.485 ;
        RECT 2.245 0.255 2.475 0.655 ;
        RECT 2.645 0.255 3.135 0.825 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__o31a_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o31a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.370 0.995 1.760 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.990 1.325 2.190 2.125 ;
        RECT 1.945 0.995 2.190 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.390 0.995 2.640 2.125 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.855 0.995 3.255 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.550 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.577500 ;
    PORT
      LAYER li1 ;
        RECT 0.550 1.835 0.990 2.465 ;
        RECT 0.550 1.295 0.860 1.835 ;
        RECT 0.085 1.075 0.860 1.295 ;
        RECT 0.550 0.825 0.860 1.075 ;
        RECT 0.550 0.265 0.990 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.465 0.380 2.635 ;
        RECT 1.165 1.785 1.480 2.635 ;
        RECT 1.650 2.295 3.080 2.465 ;
        RECT 1.650 1.615 1.820 2.295 ;
        RECT 1.030 1.445 1.820 1.615 ;
        RECT 2.830 1.665 3.080 2.295 ;
        RECT 3.255 1.835 3.590 2.635 ;
        RECT 2.830 1.495 3.595 1.665 ;
        RECT 1.030 0.995 1.200 1.445 ;
        RECT 0.085 0.085 0.380 0.905 ;
        RECT 3.425 0.825 3.595 1.495 ;
        RECT 1.160 0.085 1.610 0.825 ;
        RECT 1.780 0.655 2.940 0.825 ;
        RECT 1.780 0.255 1.950 0.655 ;
        RECT 2.120 0.085 2.540 0.485 ;
        RECT 2.710 0.255 2.940 0.655 ;
        RECT 3.110 0.255 3.595 0.825 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__o31a_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o31a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 5.140 1.055 5.470 1.360 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.680 1.530 6.355 1.700 ;
        RECT 4.680 1.360 4.970 1.530 ;
        RECT 4.265 1.055 4.970 1.360 ;
        RECT 5.640 1.055 6.355 1.530 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.765 1.055 4.095 1.360 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.780 1.355 3.150 1.695 ;
        RECT 2.780 1.055 3.575 1.355 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.120 0.105 6.280 1.015 ;
        RECT 0.125 -0.085 0.295 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.680 1.665 0.895 2.465 ;
        RECT 1.565 1.665 1.750 2.465 ;
        RECT 0.085 1.460 1.750 1.665 ;
        RECT 0.085 0.885 0.735 1.460 ;
        RECT 0.085 0.715 1.765 0.885 ;
        RECT 0.680 0.655 1.765 0.715 ;
        RECT 0.680 0.255 0.895 0.655 ;
        RECT 1.565 0.255 1.765 0.655 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.085 1.835 0.510 2.635 ;
        RECT 1.065 1.835 1.395 2.635 ;
        RECT 1.920 1.460 2.250 2.635 ;
        RECT 2.440 2.070 2.610 2.465 ;
        RECT 2.780 2.240 3.110 2.635 ;
        RECT 3.760 2.070 4.090 2.465 ;
        RECT 2.440 1.870 4.090 2.070 ;
        RECT 2.440 1.290 2.610 1.870 ;
        RECT 4.260 1.700 4.510 2.465 ;
        RECT 4.680 2.070 4.850 2.465 ;
        RECT 5.020 2.240 5.350 2.635 ;
        RECT 5.520 2.070 5.720 2.465 ;
        RECT 4.680 1.870 5.720 2.070 ;
        RECT 5.890 1.870 6.355 2.465 ;
        RECT 3.320 1.530 4.510 1.700 ;
        RECT 0.905 1.055 2.610 1.290 ;
        RECT 2.440 0.885 2.610 1.055 ;
        RECT 0.085 0.085 0.510 0.545 ;
        RECT 1.065 0.085 1.395 0.485 ;
        RECT 1.935 0.085 2.250 0.885 ;
        RECT 2.440 0.635 3.210 0.885 ;
        RECT 3.380 0.635 6.355 0.885 ;
        RECT 3.380 0.465 3.570 0.635 ;
        RECT 2.440 0.255 3.570 0.465 ;
        RECT 3.760 0.085 4.090 0.445 ;
        RECT 4.260 0.255 4.430 0.635 ;
        RECT 4.600 0.085 4.930 0.445 ;
        RECT 5.100 0.255 5.270 0.635 ;
        RECT 5.440 0.085 5.770 0.445 ;
        RECT 5.940 0.255 6.355 0.635 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 4.285 2.125 4.455 2.295 ;
        RECT 6.125 2.125 6.295 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
      LAYER met1 ;
        RECT 4.225 2.280 4.515 2.325 ;
        RECT 6.065 2.280 6.355 2.325 ;
        RECT 4.225 2.140 6.355 2.280 ;
        RECT 4.225 2.095 4.515 2.140 ;
        RECT 6.065 2.095 6.355 2.140 ;
  END
END sky130_fd_sc_hd__o31a_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o31ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.440 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.610 1.075 1.055 2.465 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.460 1.325 1.700 2.405 ;
        RECT 1.225 1.075 1.700 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.330 0.995 2.675 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.615 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.006000 ;
    PORT
      LAYER li1 ;
        RECT 1.945 0.825 2.160 2.465 ;
        RECT 1.945 0.260 2.675 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.090 1.495 0.440 2.635 ;
        RECT 2.330 1.495 2.675 2.635 ;
        RECT 0.175 0.085 0.345 0.905 ;
        RECT 0.515 0.735 1.700 0.905 ;
        RECT 0.515 0.255 0.845 0.735 ;
        RECT 1.015 0.085 1.185 0.565 ;
        RECT 1.370 0.255 1.700 0.735 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__o31ai_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o31ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.055 1.240 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.410 1.055 2.220 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.390 1.055 3.205 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.175 0.755 4.515 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.555 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.063500 ;
    PORT
      LAYER li1 ;
        RECT 2.335 1.665 2.665 2.125 ;
        RECT 3.175 1.665 3.505 2.465 ;
        RECT 4.175 1.665 4.515 2.465 ;
        RECT 2.335 1.495 4.515 1.665 ;
        RECT 3.675 0.595 4.005 1.495 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.090 1.665 0.445 2.465 ;
        RECT 0.615 1.835 0.785 2.635 ;
        RECT 0.955 1.665 1.285 2.465 ;
        RECT 1.455 2.295 3.005 2.465 ;
        RECT 1.455 1.835 1.625 2.295 ;
        RECT 1.795 1.665 2.125 2.125 ;
        RECT 2.835 1.835 3.005 2.295 ;
        RECT 3.675 1.835 4.005 2.635 ;
        RECT 0.090 1.495 2.125 1.665 ;
        RECT 0.090 0.715 3.505 0.885 ;
        RECT 0.090 0.255 0.445 0.715 ;
        RECT 0.615 0.085 0.785 0.545 ;
        RECT 0.955 0.255 1.285 0.715 ;
        RECT 1.455 0.085 1.965 0.545 ;
        RECT 2.175 0.255 2.505 0.715 ;
        RECT 2.675 0.085 3.005 0.545 ;
        RECT 3.175 0.425 3.505 0.715 ;
        RECT 4.175 0.425 4.515 0.585 ;
        RECT 3.175 0.255 4.515 0.425 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__o31ai_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o31ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o31ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.055 1.780 1.425 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.950 1.055 3.605 1.425 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.775 1.055 5.940 1.275 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.465 1.055 7.735 1.275 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.025 0.105 7.790 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.683800 ;
    PORT
      LAYER li1 ;
        RECT 5.770 1.695 5.940 2.465 ;
        RECT 6.610 1.695 6.780 2.465 ;
        RECT 7.450 1.695 7.735 2.465 ;
        RECT 3.775 1.445 7.735 1.695 ;
        RECT 6.110 0.885 6.295 1.445 ;
        RECT 6.110 0.645 7.280 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.090 1.895 0.445 2.465 ;
        RECT 0.615 2.065 0.785 2.635 ;
        RECT 0.955 1.895 1.285 2.465 ;
        RECT 1.455 2.065 1.625 2.635 ;
        RECT 1.795 2.205 3.885 2.465 ;
        RECT 1.795 1.895 2.125 2.205 ;
        RECT 0.090 1.595 2.125 1.895 ;
        RECT 2.295 1.765 2.465 2.035 ;
        RECT 2.635 1.935 2.965 2.205 ;
        RECT 4.080 2.035 5.600 2.465 ;
        RECT 3.135 1.865 5.600 2.035 ;
        RECT 6.110 1.890 6.440 2.635 ;
        RECT 6.950 1.890 7.280 2.635 ;
        RECT 3.135 1.765 3.605 1.865 ;
        RECT 2.295 1.595 3.605 1.765 ;
        RECT 0.090 0.715 5.940 0.885 ;
        RECT 0.090 0.255 0.445 0.715 ;
        RECT 0.615 0.085 0.785 0.545 ;
        RECT 0.955 0.255 1.285 0.715 ;
        RECT 1.455 0.085 1.625 0.545 ;
        RECT 1.795 0.255 2.125 0.715 ;
        RECT 2.295 0.085 2.465 0.545 ;
        RECT 2.635 0.255 2.965 0.715 ;
        RECT 3.135 0.085 3.305 0.545 ;
        RECT 3.475 0.255 3.805 0.715 ;
        RECT 3.995 0.085 4.640 0.545 ;
        RECT 4.810 0.395 4.980 0.715 ;
        RECT 5.150 0.085 5.600 0.545 ;
        RECT 5.770 0.475 5.940 0.715 ;
        RECT 7.450 0.475 7.735 0.885 ;
        RECT 5.770 0.255 7.735 0.475 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
  END
END sky130_fd_sc_hd__o31ai_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o32a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.005 1.075 1.255 1.325 ;
        RECT 1.005 0.995 1.175 1.075 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.485 1.325 1.810 2.125 ;
        RECT 1.465 0.995 1.810 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.980 0.995 2.255 1.660 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.320 0.995 3.595 1.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.440 0.995 2.795 1.660 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.175 0.105 3.675 1.015 ;
        RECT 0.175 0.085 0.310 0.105 ;
        RECT 0.140 -0.085 0.310 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.504000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.495 0.470 2.455 ;
        RECT 0.085 0.825 0.260 1.495 ;
        RECT 0.085 0.255 0.595 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.685 1.835 0.975 2.635 ;
        RECT 1.145 2.295 2.510 2.465 ;
        RECT 1.145 1.665 1.315 2.295 ;
        RECT 2.180 2.085 2.510 2.295 ;
        RECT 2.180 1.835 3.135 2.085 ;
        RECT 0.640 1.495 1.315 1.665 ;
        RECT 0.640 1.325 0.810 1.495 ;
        RECT 0.445 1.075 0.810 1.325 ;
        RECT 0.445 0.995 0.635 1.075 ;
        RECT 2.965 0.825 3.135 1.835 ;
        RECT 3.305 1.495 3.595 2.635 ;
        RECT 1.140 0.655 2.540 0.825 ;
        RECT 0.765 0.085 0.935 0.645 ;
        RECT 1.140 0.255 1.470 0.655 ;
        RECT 1.645 0.085 1.975 0.485 ;
        RECT 2.210 0.465 2.540 0.655 ;
        RECT 2.710 0.635 3.135 0.825 ;
        RECT 3.305 0.465 3.595 0.735 ;
        RECT 2.210 0.255 3.595 0.465 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__o32a_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o32a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.495 0.995 1.715 1.615 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.995 2.160 1.615 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.415 0.995 2.635 1.615 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.725 1.245 4.055 1.325 ;
        RECT 3.695 1.075 4.055 1.245 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.910 0.995 3.155 1.615 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.135 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.845 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 1.015 2.125 1.525 2.635 ;
        RECT 2.695 1.955 3.025 2.465 ;
        RECT 1.015 1.785 3.525 1.955 ;
        RECT 1.015 0.995 1.325 1.785 ;
        RECT 0.085 0.085 0.345 0.885 ;
        RECT 3.325 0.825 3.525 1.785 ;
        RECT 3.695 1.495 4.055 2.635 ;
        RECT 1.095 0.085 1.425 0.825 ;
        RECT 1.695 0.655 3.025 0.825 ;
        RECT 1.695 0.255 2.025 0.655 ;
        RECT 2.195 0.085 2.525 0.485 ;
        RECT 2.695 0.425 3.025 0.655 ;
        RECT 3.195 0.595 3.525 0.825 ;
        RECT 3.695 0.425 4.055 0.905 ;
        RECT 2.695 0.255 4.055 0.425 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__o32a_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o32a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.150 1.075 0.780 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.070 1.075 1.700 1.275 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.010 1.075 2.625 1.275 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.870 1.075 4.230 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.790 1.075 5.260 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.985 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 6.305 1.665 6.635 2.465 ;
        RECT 7.145 1.665 7.475 2.465 ;
        RECT 6.305 1.495 8.135 1.665 ;
        RECT 7.645 0.905 8.135 1.495 ;
        RECT 6.305 0.715 8.135 0.905 ;
        RECT 6.305 0.255 6.635 0.715 ;
        RECT 7.145 0.255 7.475 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.085 1.665 0.425 2.465 ;
        RECT 0.595 1.835 0.765 2.635 ;
        RECT 0.935 2.295 2.105 2.465 ;
        RECT 0.935 1.665 1.265 2.295 ;
        RECT 0.085 1.445 1.265 1.665 ;
        RECT 1.435 1.690 1.605 2.045 ;
        RECT 1.775 1.860 2.105 2.295 ;
        RECT 2.295 2.295 3.465 2.465 ;
        RECT 2.295 1.690 2.625 2.295 ;
        RECT 1.435 1.445 2.625 1.690 ;
        RECT 2.795 1.275 2.965 2.045 ;
        RECT 3.135 1.445 3.465 2.295 ;
        RECT 3.655 1.955 3.985 2.465 ;
        RECT 4.155 2.125 4.325 2.635 ;
        RECT 4.495 2.285 5.695 2.465 ;
        RECT 4.495 1.955 4.825 2.285 ;
        RECT 3.655 1.785 4.825 1.955 ;
        RECT 3.655 1.445 3.985 1.785 ;
        RECT 5.025 1.615 5.195 2.115 ;
        RECT 4.400 1.445 5.195 1.615 ;
        RECT 5.365 1.445 5.695 2.285 ;
        RECT 5.965 1.835 6.135 2.635 ;
        RECT 6.805 1.835 6.975 2.635 ;
        RECT 7.645 1.835 7.900 2.635 ;
        RECT 2.795 1.105 3.645 1.275 ;
        RECT 0.085 0.635 2.965 0.885 ;
        RECT 3.455 0.805 3.645 1.105 ;
        RECT 4.400 0.805 4.620 1.445 ;
        RECT 5.520 1.245 6.135 1.265 ;
        RECT 5.520 1.075 7.475 1.245 ;
        RECT 5.520 0.805 5.775 1.075 ;
        RECT 3.455 0.635 5.775 0.805 ;
        RECT 0.085 0.255 0.345 0.635 ;
        RECT 2.715 0.465 2.965 0.635 ;
        RECT 0.515 0.085 2.545 0.465 ;
        RECT 2.715 0.255 5.695 0.465 ;
        RECT 5.965 0.085 6.135 0.885 ;
        RECT 6.805 0.085 6.975 0.545 ;
        RECT 7.645 0.085 7.900 0.545 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
  END
END sky130_fd_sc_hd__o32a_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o32ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.575 0.995 3.135 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.930 0.995 2.225 2.465 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.410 0.995 1.700 1.615 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.995 0.360 1.325 ;
        RECT 0.090 0.685 0.345 0.995 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.870 0.995 1.240 1.615 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.215 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.821250 ;
    PORT
      LAYER li1 ;
        RECT 0.530 1.785 1.545 2.465 ;
        RECT 0.530 0.825 0.700 1.785 ;
        RECT 0.515 0.655 0.845 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.090 1.495 0.360 2.635 ;
        RECT 2.695 1.495 3.135 2.635 ;
        RECT 1.015 0.655 2.525 0.825 ;
        RECT 1.015 0.485 1.345 0.655 ;
        RECT 0.090 0.255 1.345 0.485 ;
        RECT 1.515 0.085 2.185 0.485 ;
        RECT 2.355 0.375 2.525 0.655 ;
        RECT 2.695 0.085 3.135 0.825 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__o32ai_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o32ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.750 1.075 5.865 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.370 1.075 4.480 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.075 3.065 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.075 1.705 1.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.845 1.325 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.845 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.095 ;
        RECT 2.775 1.665 3.105 2.085 ;
        RECT 0.515 1.495 3.105 1.665 ;
        RECT 1.875 1.105 2.170 1.495 ;
        RECT 1.875 0.905 2.045 1.105 ;
        RECT 0.515 0.655 2.045 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.090 2.295 1.265 2.465 ;
        RECT 0.090 1.495 0.345 2.295 ;
        RECT 1.015 2.005 1.265 2.295 ;
        RECT 1.435 2.175 1.605 2.635 ;
        RECT 1.775 2.005 2.105 2.455 ;
        RECT 1.015 1.835 2.105 2.005 ;
        RECT 2.335 2.255 4.385 2.445 ;
        RECT 2.335 1.835 2.585 2.255 ;
        RECT 3.275 1.495 3.445 2.255 ;
        RECT 3.615 1.665 3.945 2.085 ;
        RECT 4.135 1.835 4.385 2.255 ;
        RECT 4.620 1.835 4.825 2.635 ;
        RECT 4.995 1.665 5.325 2.460 ;
        RECT 3.615 1.495 5.325 1.665 ;
        RECT 5.495 1.495 5.715 2.635 ;
        RECT 0.090 0.485 0.345 0.905 ;
        RECT 2.235 0.715 5.755 0.905 ;
        RECT 2.235 0.485 2.405 0.715 ;
        RECT 0.090 0.255 2.405 0.485 ;
        RECT 2.620 0.085 2.950 0.545 ;
        RECT 3.135 0.255 3.465 0.715 ;
        RECT 3.635 0.085 3.805 0.545 ;
        RECT 4.055 0.255 4.725 0.715 ;
        RECT 4.905 0.085 5.235 0.545 ;
        RECT 5.425 0.255 5.755 0.715 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
END sky130_fd_sc_hd__o32ai_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o32ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o32ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 8.290 1.075 10.035 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.090 1.075 7.260 1.275 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.770 1.075 5.380 1.275 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 2.205 1.075 3.540 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.110 1.075 1.685 1.275 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 10.065 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.085 ;
        RECT 1.355 1.665 1.700 2.085 ;
        RECT 4.410 1.665 4.740 2.085 ;
        RECT 5.250 1.665 5.580 2.085 ;
        RECT 0.515 1.495 5.580 1.665 ;
        RECT 1.855 0.905 2.035 1.495 ;
        RECT 0.515 0.655 3.380 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.090 2.255 2.040 2.465 ;
        RECT 0.090 1.495 0.345 2.255 ;
        RECT 1.015 1.835 1.185 2.255 ;
        RECT 1.870 2.005 2.040 2.255 ;
        RECT 2.210 2.175 2.540 2.635 ;
        RECT 2.710 2.005 2.880 2.425 ;
        RECT 3.050 2.175 3.380 2.635 ;
        RECT 3.550 2.005 3.800 2.465 ;
        RECT 1.870 1.835 3.800 2.005 ;
        RECT 3.990 2.255 7.680 2.465 ;
        RECT 3.990 1.835 4.240 2.255 ;
        RECT 4.910 1.835 5.080 2.255 ;
        RECT 5.750 1.835 5.920 2.255 ;
        RECT 6.090 1.665 6.420 2.085 ;
        RECT 6.590 1.835 6.760 2.255 ;
        RECT 6.930 1.665 7.260 2.085 ;
        RECT 7.430 1.835 7.680 2.255 ;
        RECT 7.870 1.835 8.120 2.635 ;
        RECT 8.290 1.665 8.620 2.465 ;
        RECT 8.790 1.835 8.960 2.635 ;
        RECT 9.130 1.665 9.460 2.465 ;
        RECT 6.090 1.495 9.460 1.665 ;
        RECT 9.630 1.495 10.035 2.635 ;
        RECT 0.090 0.465 0.345 0.905 ;
        RECT 3.550 0.735 10.035 0.905 ;
        RECT 3.550 0.465 3.800 0.735 ;
        RECT 0.090 0.255 3.800 0.465 ;
        RECT 3.970 0.085 4.140 0.545 ;
        RECT 4.310 0.255 4.640 0.735 ;
        RECT 4.810 0.085 5.140 0.545 ;
        RECT 5.310 0.255 5.980 0.735 ;
        RECT 6.170 0.085 6.340 0.545 ;
        RECT 6.510 0.255 6.840 0.735 ;
        RECT 7.010 0.085 7.180 0.545 ;
        RECT 7.350 0.255 8.040 0.735 ;
        RECT 8.370 0.085 8.540 0.545 ;
        RECT 8.710 0.255 9.040 0.735 ;
        RECT 9.210 0.085 9.470 0.545 ;
        RECT 9.645 0.255 10.035 0.735 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
  END
END sky130_fd_sc_hd__o32ai_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o41a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.485 1.075 3.995 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.075 3.275 2.390 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.075 2.735 2.390 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.865 1.075 2.195 2.390 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.275 1.075 1.695 1.285 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.065 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.672000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.455 0.610 2.465 ;
        RECT 0.085 0.885 0.355 1.455 ;
        RECT 0.085 0.255 0.425 0.885 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.845 1.915 1.175 2.635 ;
        RECT 1.345 1.745 1.595 2.465 ;
        RECT 0.845 1.455 1.595 1.745 ;
        RECT 3.605 1.515 3.935 2.635 ;
        RECT 0.845 1.285 1.105 1.455 ;
        RECT 0.525 1.075 1.105 1.285 ;
        RECT 0.735 0.905 1.105 1.075 ;
        RECT 0.735 0.715 1.485 0.905 ;
        RECT 0.715 0.085 0.885 0.545 ;
        RECT 1.155 0.270 1.485 0.715 ;
        RECT 1.655 0.735 3.955 0.905 ;
        RECT 1.655 0.415 1.825 0.735 ;
        RECT 2.050 0.085 2.380 0.545 ;
        RECT 2.580 0.255 2.910 0.735 ;
        RECT 3.125 0.085 3.455 0.545 ;
        RECT 3.625 0.255 3.955 0.735 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__o41a_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o41a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.825 1.075 4.515 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.325 1.075 3.655 2.335 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.825 1.075 3.155 2.340 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.075 2.655 2.340 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.775 1.075 2.155 1.325 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.525 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.495 0.845 2.465 ;
        RECT 0.515 0.880 0.790 1.495 ;
        RECT 0.515 0.255 0.845 0.880 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.525 2.635 ;
        RECT 1.015 1.495 1.185 1.835 ;
        RECT 1.695 1.665 2.145 2.465 ;
        RECT 1.355 1.495 2.145 1.665 ;
        RECT 4.065 1.495 4.395 2.635 ;
        RECT 1.355 1.325 1.600 1.495 ;
        RECT 0.960 1.075 1.600 1.325 ;
        RECT 0.085 0.085 0.345 0.885 ;
        RECT 1.015 0.085 1.260 0.885 ;
        RECT 1.430 0.850 1.600 1.075 ;
        RECT 1.430 0.255 1.785 0.850 ;
        RECT 1.985 0.715 4.395 0.905 ;
        RECT 1.985 0.255 2.315 0.715 ;
        RECT 2.485 0.085 2.750 0.545 ;
        RECT 2.955 0.255 3.285 0.715 ;
        RECT 3.505 0.085 3.775 0.545 ;
        RECT 4.065 0.255 4.395 0.715 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__o41a_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o41a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 6.650 1.075 7.735 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 5.150 1.075 6.360 1.275 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.330 1.075 4.960 1.275 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.410 1.075 4.040 1.275 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.835 1.075 3.165 1.275 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.725 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.355 1.665 1.685 2.465 ;
        RECT 0.085 1.465 1.685 1.665 ;
        RECT 0.085 0.905 0.345 1.465 ;
        RECT 0.085 0.715 1.685 0.905 ;
        RECT 0.515 0.255 0.845 0.715 ;
        RECT 1.355 0.255 1.685 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.085 1.835 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.465 2.025 2.635 ;
        RECT 2.195 1.615 2.545 2.465 ;
        RECT 2.715 1.835 2.965 2.635 ;
        RECT 3.135 2.295 4.325 2.465 ;
        RECT 3.135 1.835 3.405 2.295 ;
        RECT 3.575 1.615 3.825 2.125 ;
        RECT 2.195 1.445 3.825 1.615 ;
        RECT 3.995 1.615 4.325 2.295 ;
        RECT 4.495 2.295 6.145 2.465 ;
        RECT 4.495 1.785 4.665 2.295 ;
        RECT 4.835 1.615 5.165 2.115 ;
        RECT 3.995 1.445 5.165 1.615 ;
        RECT 5.395 1.615 5.645 2.115 ;
        RECT 5.815 1.785 6.145 2.295 ;
        RECT 6.315 1.615 6.485 2.455 ;
        RECT 6.655 1.785 6.985 2.635 ;
        RECT 7.265 1.615 7.595 2.465 ;
        RECT 5.395 1.445 7.595 1.615 ;
        RECT 2.195 1.295 2.545 1.445 ;
        RECT 0.515 1.245 2.545 1.295 ;
        RECT 0.515 1.075 2.665 1.245 ;
        RECT 2.295 0.905 2.665 1.075 ;
        RECT 0.085 0.085 0.345 0.545 ;
        RECT 1.015 0.085 1.185 0.545 ;
        RECT 1.855 0.085 2.105 0.885 ;
        RECT 2.295 0.635 3.045 0.905 ;
        RECT 3.235 0.735 7.595 0.905 ;
        RECT 3.235 0.465 3.485 0.735 ;
        RECT 2.295 0.255 3.485 0.465 ;
        RECT 3.655 0.085 3.875 0.545 ;
        RECT 4.075 0.255 4.245 0.735 ;
        RECT 4.445 0.085 4.715 0.545 ;
        RECT 4.915 0.255 5.085 0.735 ;
        RECT 5.305 0.085 5.915 0.545 ;
        RECT 6.240 0.255 6.410 0.735 ;
        RECT 6.685 0.085 6.955 0.545 ;
        RECT 7.265 0.255 7.595 0.735 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
  END
END sky130_fd_sc_hd__o41a_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o41ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.500 1.075 3.080 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.990 1.415 2.330 2.355 ;
        RECT 2.000 1.075 2.330 1.415 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.500 1.245 1.820 2.355 ;
        RECT 1.500 1.075 1.830 1.245 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.015 1.245 1.320 2.355 ;
        RECT 0.990 1.075 1.320 1.245 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.440 1.275 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.070 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.439000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.485 0.845 2.465 ;
        RECT 0.610 0.905 0.780 1.485 ;
        RECT 0.085 0.735 0.780 0.905 ;
        RECT 0.085 0.255 0.425 0.735 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.445 0.345 2.635 ;
        RECT 2.630 1.495 2.960 2.635 ;
        RECT 0.950 0.735 2.960 0.905 ;
        RECT 0.950 0.565 1.120 0.735 ;
        RECT 0.790 0.255 1.120 0.565 ;
        RECT 1.290 0.085 1.540 0.565 ;
        RECT 1.710 0.255 2.040 0.735 ;
        RECT 2.210 0.085 2.460 0.565 ;
        RECT 2.630 0.255 2.960 0.735 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__o41ai_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o41ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.720 1.075 5.895 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.780 1.075 4.540 1.275 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.595 1.075 3.580 1.275 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.500 1.075 2.325 1.275 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 0.440 1.275 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.815 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.715500 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.665 0.845 2.465 ;
        RECT 1.875 1.665 2.205 2.125 ;
        RECT 0.515 1.505 2.205 1.665 ;
        RECT 0.610 1.445 2.205 1.505 ;
        RECT 0.610 0.885 0.845 1.445 ;
        RECT 0.515 0.635 0.845 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 1.015 1.835 1.265 2.635 ;
        RECT 1.455 2.295 2.545 2.465 ;
        RECT 1.455 1.835 1.705 2.295 ;
        RECT 2.375 1.615 2.545 2.295 ;
        RECT 2.715 2.295 4.445 2.465 ;
        RECT 2.715 1.835 3.045 2.295 ;
        RECT 3.215 1.615 3.465 2.125 ;
        RECT 2.375 1.445 3.465 1.615 ;
        RECT 3.695 1.615 3.945 2.125 ;
        RECT 4.115 1.835 4.445 2.295 ;
        RECT 4.615 1.615 4.785 2.465 ;
        RECT 4.955 1.785 5.285 2.635 ;
        RECT 5.455 1.615 5.705 2.465 ;
        RECT 3.695 1.445 5.705 1.615 ;
        RECT 0.085 0.465 0.345 0.905 ;
        RECT 1.015 0.735 5.705 0.905 ;
        RECT 1.015 0.465 1.265 0.735 ;
        RECT 0.085 0.255 1.265 0.465 ;
        RECT 1.455 0.085 1.705 0.545 ;
        RECT 1.875 0.255 2.205 0.735 ;
        RECT 2.375 0.085 2.545 0.545 ;
        RECT 2.715 0.255 3.045 0.735 ;
        RECT 3.215 0.085 3.450 0.545 ;
        RECT 3.695 0.255 4.025 0.735 ;
        RECT 4.195 0.085 4.365 0.545 ;
        RECT 4.535 0.255 4.865 0.735 ;
        RECT 5.035 0.085 5.205 0.545 ;
        RECT 5.375 0.255 5.705 0.735 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
END sky130_fd_sc_hd__o41ai_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o41ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o41ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 8.155 1.075 10.035 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.170 1.075 7.940 1.275 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 4.310 1.075 5.980 1.275 ;
    END
  END A3
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 2.350 1.075 4.020 1.275 ;
    END
  END A4
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 1.075 1.700 1.275 ;
    END
  END B1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.975 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.431000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 1.615 0.845 2.465 ;
        RECT 1.355 1.615 1.685 2.465 ;
        RECT 2.715 1.615 3.045 2.125 ;
        RECT 3.555 1.615 3.885 2.125 ;
        RECT 0.515 1.445 3.885 1.615 ;
        RECT 1.870 0.905 2.160 1.445 ;
        RECT 0.515 0.635 2.160 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.085 1.445 0.345 2.635 ;
        RECT 1.015 1.835 1.185 2.635 ;
        RECT 1.855 1.835 2.105 2.635 ;
        RECT 2.295 2.295 4.225 2.465 ;
        RECT 2.295 1.785 2.545 2.295 ;
        RECT 3.215 1.785 3.385 2.295 ;
        RECT 4.055 1.615 4.225 2.295 ;
        RECT 4.395 2.295 7.685 2.465 ;
        RECT 4.395 1.785 4.645 2.295 ;
        RECT 4.815 1.615 5.145 2.125 ;
        RECT 5.315 1.785 5.485 2.295 ;
        RECT 5.655 1.615 5.985 2.125 ;
        RECT 4.055 1.445 5.985 1.615 ;
        RECT 6.175 1.615 6.505 2.125 ;
        RECT 6.675 1.785 6.845 2.295 ;
        RECT 7.015 1.615 7.345 2.125 ;
        RECT 7.515 1.785 7.685 2.295 ;
        RECT 7.855 1.615 8.185 2.465 ;
        RECT 8.355 1.835 8.525 2.635 ;
        RECT 8.695 1.615 9.025 2.465 ;
        RECT 9.195 1.835 9.365 2.635 ;
        RECT 9.535 1.615 9.865 2.465 ;
        RECT 6.175 1.445 9.865 1.615 ;
        RECT 0.085 0.465 0.345 0.905 ;
        RECT 2.350 0.735 9.865 0.905 ;
        RECT 2.350 0.465 2.625 0.735 ;
        RECT 0.085 0.255 2.625 0.465 ;
        RECT 2.795 0.085 2.965 0.545 ;
        RECT 3.135 0.255 3.465 0.735 ;
        RECT 3.635 0.085 3.805 0.545 ;
        RECT 3.975 0.255 4.305 0.735 ;
        RECT 4.475 0.085 4.645 0.545 ;
        RECT 4.815 0.255 5.145 0.735 ;
        RECT 5.315 0.085 5.485 0.545 ;
        RECT 5.655 0.255 5.985 0.735 ;
        RECT 6.175 0.260 6.505 0.735 ;
        RECT 6.675 0.085 6.845 0.545 ;
        RECT 7.015 0.260 7.345 0.735 ;
        RECT 7.515 0.085 7.685 0.545 ;
        RECT 7.855 0.260 8.185 0.735 ;
        RECT 8.355 0.085 8.525 0.545 ;
        RECT 8.695 0.260 9.025 0.735 ;
        RECT 9.195 0.085 9.365 0.545 ;
        RECT 9.535 0.260 9.865 0.735 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
  END
END sky130_fd_sc_hd__o41ai_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o211a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.300 1.075 1.720 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.890 1.075 2.220 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.390 1.075 2.720 1.275 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.245 1.075 3.595 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.480 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.495 0.425 2.465 ;
        RECT 0.085 0.885 0.260 1.495 ;
        RECT 0.085 0.255 0.425 0.885 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.595 1.495 0.765 2.635 ;
        RECT 1.035 1.835 1.285 2.635 ;
        RECT 1.930 1.665 2.260 2.465 ;
        RECT 2.560 1.835 2.890 2.635 ;
        RECT 3.060 1.665 3.390 2.465 ;
        RECT 0.955 1.495 3.390 1.665 ;
        RECT 0.955 1.245 1.125 1.495 ;
        RECT 0.430 1.075 1.125 1.245 ;
        RECT 0.595 0.085 0.845 0.885 ;
        RECT 1.035 0.735 2.260 0.905 ;
        RECT 1.035 0.255 1.365 0.735 ;
        RECT 1.535 0.085 1.760 0.545 ;
        RECT 1.930 0.255 2.260 0.735 ;
        RECT 2.890 0.865 3.060 1.495 ;
        RECT 2.890 0.255 3.390 0.865 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__o211a_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o211a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.990 0.995 2.325 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.530 0.995 1.820 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.880 0.995 1.240 1.325 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.360 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.660 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER li1 ;
        RECT 2.810 2.075 3.000 2.465 ;
        RECT 2.810 1.905 3.540 2.075 ;
        RECT 3.345 0.785 3.540 1.905 ;
        RECT 2.720 0.615 3.540 0.785 ;
        RECT 2.720 0.255 3.050 0.615 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.090 1.765 0.355 2.465 ;
        RECT 0.525 1.935 0.855 2.635 ;
        RECT 1.025 1.765 1.695 2.465 ;
        RECT 2.200 1.935 2.630 2.635 ;
        RECT 3.170 2.255 3.500 2.635 ;
        RECT 0.090 1.510 2.665 1.765 ;
        RECT 0.530 0.825 0.710 1.510 ;
        RECT 2.495 1.325 2.665 1.510 ;
        RECT 2.495 0.995 3.175 1.325 ;
        RECT 0.095 0.425 0.710 0.825 ;
        RECT 0.880 0.635 2.150 0.825 ;
        RECT 0.095 0.255 0.430 0.425 ;
        RECT 1.390 0.085 1.725 0.465 ;
        RECT 2.315 0.085 2.550 0.525 ;
        RECT 3.220 0.085 3.550 0.445 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__o211a_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o211a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.490 1.495 6.290 1.685 ;
        RECT 4.490 1.035 4.845 1.495 ;
        RECT 5.890 1.035 6.290 1.495 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 5.030 1.035 5.705 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.540 1.445 4.280 1.685 ;
        RECT 2.540 0.995 2.830 1.445 ;
        RECT 3.950 1.035 4.280 1.445 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.055 1.035 3.740 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.435 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.630 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.911000 ;
    PORT
      LAYER li1 ;
        RECT 0.980 1.700 1.160 2.465 ;
        RECT 1.840 1.700 2.030 2.465 ;
        RECT 0.085 1.435 2.030 1.700 ;
        RECT 0.085 0.805 0.365 1.435 ;
        RECT 0.085 0.635 1.605 0.805 ;
        RECT 0.595 0.615 1.605 0.635 ;
        RECT 0.595 0.255 0.765 0.615 ;
        RECT 1.435 0.255 1.605 0.615 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.440 2.805 ;
        RECT 0.480 1.870 0.810 2.635 ;
        RECT 1.340 1.870 1.670 2.635 ;
        RECT 2.200 2.200 2.530 2.635 ;
        RECT 2.700 2.025 3.060 2.465 ;
        RECT 3.285 2.195 3.615 2.635 ;
        RECT 3.785 2.025 4.120 2.465 ;
        RECT 4.290 2.195 4.555 2.635 ;
        RECT 5.155 2.025 5.485 2.465 ;
        RECT 2.200 1.855 5.485 2.025 ;
        RECT 6.015 1.915 6.345 2.635 ;
        RECT 2.200 1.265 2.370 1.855 ;
        RECT 0.535 1.065 2.370 1.265 ;
        RECT 2.200 0.815 2.370 1.065 ;
        RECT 2.200 0.635 3.520 0.815 ;
        RECT 4.170 0.695 6.345 0.865 ;
        RECT 4.170 0.465 4.500 0.695 ;
        RECT 0.095 0.085 0.425 0.465 ;
        RECT 0.935 0.085 1.265 0.445 ;
        RECT 1.775 0.085 2.140 0.465 ;
        RECT 2.330 0.255 4.500 0.465 ;
        RECT 4.670 0.085 4.985 0.525 ;
        RECT 5.155 0.255 5.485 0.695 ;
        RECT 5.655 0.085 5.845 0.525 ;
        RECT 6.015 0.255 6.345 0.695 ;
        RECT 0.000 -0.085 6.440 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
  END
END sky130_fd_sc_hd__o211a_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o211ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.395 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.325 0.775 2.250 ;
        RECT 0.605 0.995 0.980 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.470 1.325 1.795 1.615 ;
        RECT 1.300 0.995 1.795 1.325 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.970 1.075 2.300 1.615 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 2.725 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.418250 ;
    PORT
      LAYER li1 ;
        RECT 0.945 2.045 1.275 2.445 ;
        RECT 1.975 2.045 2.675 2.465 ;
        RECT 0.945 1.815 2.675 2.045 ;
        RECT 0.945 1.595 1.275 1.815 ;
        RECT 2.470 0.845 2.675 1.815 ;
        RECT 1.965 0.255 2.675 0.845 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.095 1.575 0.425 2.635 ;
        RECT 1.445 2.275 1.775 2.635 ;
        RECT 0.095 0.615 1.455 0.825 ;
        RECT 0.095 0.255 0.425 0.615 ;
        RECT 0.595 0.085 0.925 0.445 ;
        RECT 1.125 0.255 1.455 0.615 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__o211ai_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o211ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.560 1.245 4.455 1.295 ;
        RECT 3.505 1.075 4.455 1.245 ;
        RECT 4.115 0.765 4.455 1.075 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.365 1.075 3.335 1.355 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.075 1.905 1.365 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.375 1.970 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.555 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.022000 ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.710 0.805 2.465 ;
        RECT 1.475 1.710 1.665 2.465 ;
        RECT 2.825 1.710 3.155 2.125 ;
        RECT 0.545 1.540 3.155 1.710 ;
        RECT 0.545 0.670 0.875 1.540 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.115 2.175 0.375 2.635 ;
        RECT 0.975 1.915 1.305 2.635 ;
        RECT 1.835 1.915 2.165 2.635 ;
        RECT 2.395 2.295 3.515 2.465 ;
        RECT 2.395 2.100 2.655 2.295 ;
        RECT 3.325 1.695 3.515 2.295 ;
        RECT 3.685 1.865 4.015 2.635 ;
        RECT 4.185 1.695 4.445 2.465 ;
        RECT 3.325 1.525 4.445 1.695 ;
        RECT 1.045 0.465 1.235 0.890 ;
        RECT 1.405 0.635 3.945 0.845 ;
        RECT 3.755 0.515 3.945 0.635 ;
        RECT 1.045 0.445 2.165 0.465 ;
        RECT 0.095 0.255 2.165 0.445 ;
        RECT 2.395 0.085 2.725 0.445 ;
        RECT 3.255 0.085 3.585 0.445 ;
        RECT 4.115 0.085 4.445 0.445 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__o211ai_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o211ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o211ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.965 1.515 3.630 1.685 ;
        RECT 0.965 1.330 1.410 1.515 ;
        RECT 0.400 1.075 1.410 1.330 ;
        RECT 3.350 0.995 3.630 1.515 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.705 1.075 3.180 1.345 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 4.260 1.515 7.000 1.685 ;
        RECT 4.260 1.410 4.975 1.515 ;
        RECT 3.800 0.995 4.975 1.410 ;
        RECT 6.830 0.995 7.000 1.515 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 5.370 1.075 6.440 1.345 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.565 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.001000 ;
    PORT
      LAYER li1 ;
        RECT 1.805 2.025 3.470 2.105 ;
        RECT 4.045 2.025 7.680 2.105 ;
        RECT 1.805 1.855 7.680 2.025 ;
        RECT 7.170 1.340 7.680 1.855 ;
        RECT 7.170 0.825 7.350 1.340 ;
        RECT 6.565 0.655 7.350 0.825 ;
        RECT 6.565 0.450 6.735 0.655 ;
        RECT 5.280 0.270 6.735 0.450 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.090 1.665 0.385 2.635 ;
        RECT 0.955 2.275 1.285 2.635 ;
        RECT 1.455 2.275 3.435 2.465 ;
        RECT 0.555 2.105 0.775 2.190 ;
        RECT 1.455 2.105 1.635 2.275 ;
        RECT 3.615 2.195 3.885 2.635 ;
        RECT 4.435 2.275 4.765 2.635 ;
        RECT 5.280 2.275 5.610 2.635 ;
        RECT 6.120 2.275 6.455 2.635 ;
        RECT 7.355 2.275 7.685 2.635 ;
        RECT 0.555 1.935 1.635 2.105 ;
        RECT 0.555 1.860 0.775 1.935 ;
        RECT 0.155 0.865 1.795 0.905 ;
        RECT 0.155 0.795 3.130 0.865 ;
        RECT 0.155 0.695 3.835 0.795 ;
        RECT 0.155 0.625 1.240 0.695 ;
        RECT 1.775 0.625 3.835 0.695 ;
        RECT 4.005 0.635 6.170 0.815 ;
        RECT 0.155 0.535 0.355 0.625 ;
        RECT 0.525 0.085 0.855 0.445 ;
        RECT 1.025 0.425 1.240 0.625 ;
        RECT 1.465 0.085 1.635 0.525 ;
        RECT 3.605 0.455 3.835 0.625 ;
        RECT 7.510 0.480 7.680 0.595 ;
        RECT 2.245 0.085 2.575 0.445 ;
        RECT 3.105 0.085 3.435 0.445 ;
        RECT 3.605 0.255 4.920 0.455 ;
        RECT 6.980 0.310 7.680 0.480 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 1.070 0.425 1.240 0.595 ;
        RECT 7.510 0.425 7.680 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
      LAYER met1 ;
        RECT 1.010 0.580 1.300 0.625 ;
        RECT 7.450 0.580 7.740 0.625 ;
        RECT 1.010 0.440 7.740 0.580 ;
        RECT 1.010 0.395 1.300 0.440 ;
        RECT 7.450 0.395 7.740 0.440 ;
  END
END sky130_fd_sc_hd__o211ai_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o221a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.680 1.075 3.130 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.005 1.285 2.380 1.705 ;
        RECT 2.005 1.075 2.490 1.285 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.925 1.075 1.255 1.285 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.495 1.325 1.815 1.705 ;
        RECT 1.435 1.075 1.815 1.325 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.415 1.285 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155 0.105 3.810 1.015 ;
        RECT 0.155 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER li1 ;
        RECT 3.390 1.875 4.055 2.465 ;
        RECT 3.805 0.905 4.055 1.875 ;
        RECT 3.370 0.265 4.055 0.905 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.240 1.625 0.540 2.465 ;
        RECT 0.735 1.795 0.985 2.635 ;
        RECT 1.575 2.045 2.380 2.465 ;
        RECT 1.155 1.875 2.720 2.045 ;
        RECT 1.155 1.625 1.325 1.875 ;
        RECT 0.240 1.455 1.325 1.625 ;
        RECT 2.550 1.625 2.720 1.875 ;
        RECT 2.890 1.795 3.220 2.635 ;
        RECT 2.550 1.455 3.470 1.625 ;
        RECT 0.585 0.825 0.755 1.455 ;
        RECT 3.300 1.285 3.470 1.455 ;
        RECT 3.300 1.075 3.635 1.285 ;
        RECT 0.245 0.645 0.755 0.825 ;
        RECT 1.160 0.735 2.860 0.905 ;
        RECT 1.160 0.645 1.545 0.735 ;
        RECT 0.245 0.255 0.575 0.645 ;
        RECT 0.745 0.305 1.930 0.475 ;
        RECT 2.190 0.085 2.360 0.555 ;
        RECT 2.530 0.270 2.860 0.735 ;
        RECT 3.030 0.085 3.200 0.905 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__o221a_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o221a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.635 1.075 3.075 1.285 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.980 1.285 2.285 1.705 ;
        RECT 1.980 1.075 2.465 1.285 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.885 1.075 1.230 1.275 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.500 1.275 1.790 1.705 ;
        RECT 1.400 1.075 1.790 1.275 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.345 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.060 0.105 4.135 1.015 ;
        RECT 0.120 -0.085 0.290 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 3.295 2.045 3.545 2.465 ;
        RECT 3.295 1.875 4.055 2.045 ;
        RECT 3.745 0.905 4.055 1.875 ;
        RECT 3.295 0.735 4.055 0.905 ;
        RECT 3.295 0.265 3.625 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.250 1.670 0.580 2.465 ;
        RECT 0.750 1.850 0.990 2.635 ;
        RECT 1.550 2.045 2.305 2.465 ;
        RECT 1.160 1.875 2.625 2.045 ;
        RECT 1.160 1.670 1.330 1.875 ;
        RECT 0.250 1.495 1.330 1.670 ;
        RECT 0.545 1.445 1.330 1.495 ;
        RECT 2.455 1.625 2.625 1.875 ;
        RECT 2.795 1.795 3.125 2.635 ;
        RECT 3.715 2.215 4.055 2.635 ;
        RECT 2.455 1.455 3.415 1.625 ;
        RECT 0.545 0.805 0.715 1.445 ;
        RECT 3.245 1.285 3.415 1.455 ;
        RECT 3.245 1.075 3.575 1.285 ;
        RECT 0.170 0.635 0.715 0.805 ;
        RECT 1.085 0.735 2.785 0.905 ;
        RECT 1.085 0.645 1.470 0.735 ;
        RECT 0.170 0.255 0.500 0.635 ;
        RECT 0.670 0.295 1.855 0.465 ;
        RECT 2.115 0.085 2.285 0.555 ;
        RECT 2.455 0.270 2.785 0.735 ;
        RECT 2.955 0.085 3.125 0.905 ;
        RECT 3.795 0.085 3.965 0.565 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__o221a_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o221a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.005 1.445 4.775 1.615 ;
        RECT 3.005 1.075 3.605 1.445 ;
        RECT 4.525 1.275 4.775 1.445 ;
        RECT 4.525 1.075 5.035 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.775 1.075 4.355 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.025 1.445 2.745 1.615 ;
        RECT 1.025 1.075 1.520 1.445 ;
        RECT 2.415 1.075 2.745 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.690 1.075 2.245 1.275 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.440 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.915 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 5.315 1.955 5.525 2.465 ;
        RECT 5.315 1.785 5.900 1.955 ;
        RECT 5.730 1.615 5.900 1.785 ;
        RECT 6.115 1.615 6.365 2.465 ;
        RECT 5.730 1.445 6.920 1.615 ;
        RECT 6.575 0.905 6.920 1.445 ;
        RECT 5.235 0.735 6.920 0.905 ;
        RECT 5.235 0.725 6.405 0.735 ;
        RECT 5.235 0.255 5.565 0.725 ;
        RECT 6.075 0.255 6.405 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.145 1.455 0.395 2.635 ;
        RECT 0.565 1.955 0.815 2.465 ;
        RECT 0.985 2.125 1.235 2.635 ;
        RECT 1.405 2.295 2.495 2.465 ;
        RECT 1.405 2.125 1.655 2.295 ;
        RECT 2.245 2.125 2.495 2.295 ;
        RECT 2.665 2.125 3.425 2.635 ;
        RECT 3.595 2.295 4.685 2.465 ;
        RECT 3.595 2.125 3.845 2.295 ;
        RECT 4.435 2.125 4.685 2.295 ;
        RECT 4.855 2.125 5.105 2.635 ;
        RECT 5.695 2.125 5.945 2.635 ;
        RECT 1.825 1.955 2.075 2.125 ;
        RECT 4.015 1.955 4.265 2.125 ;
        RECT 0.565 1.785 5.145 1.955 ;
        RECT 6.535 1.795 6.785 2.635 ;
        RECT 0.565 1.445 0.845 1.785 ;
        RECT 4.975 1.615 5.145 1.785 ;
        RECT 4.975 1.445 5.375 1.615 ;
        RECT 0.085 0.475 0.345 0.895 ;
        RECT 0.610 0.865 0.845 1.445 ;
        RECT 5.205 1.275 5.375 1.445 ;
        RECT 5.205 1.075 6.405 1.275 ;
        RECT 0.515 0.645 0.845 0.865 ;
        RECT 1.015 0.475 1.185 0.905 ;
        RECT 1.355 0.725 4.725 0.905 ;
        RECT 1.355 0.715 3.885 0.725 ;
        RECT 1.355 0.645 2.535 0.715 ;
        RECT 0.085 0.255 2.955 0.475 ;
        RECT 3.145 0.085 3.385 0.545 ;
        RECT 3.555 0.255 3.885 0.715 ;
        RECT 4.055 0.085 4.225 0.555 ;
        RECT 4.395 0.255 4.725 0.725 ;
        RECT 4.895 0.085 5.065 0.905 ;
        RECT 5.735 0.085 5.905 0.555 ;
        RECT 6.575 0.085 6.830 0.565 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
END sky130_fd_sc_hd__o221a_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o221ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.675 1.075 3.135 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.465 1.615 2.675 2.405 ;
        RECT 2.295 1.445 2.675 1.615 ;
        RECT 2.295 1.245 2.505 1.445 ;
        RECT 2.165 1.075 2.505 1.245 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.010 0.995 1.355 1.325 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 1.985 1.325 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.465 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.215 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.899000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.705 0.365 2.465 ;
        RECT 1.735 1.785 2.245 2.465 ;
        RECT 1.735 1.705 2.125 1.785 ;
        RECT 0.085 1.495 2.125 1.705 ;
        RECT 0.635 0.825 0.840 1.495 ;
        RECT 0.085 0.645 0.840 0.825 ;
        RECT 0.085 0.365 0.345 0.645 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.550 1.875 1.340 2.635 ;
        RECT 2.875 1.455 3.135 2.635 ;
        RECT 2.105 0.825 3.135 0.865 ;
        RECT 1.010 0.695 3.135 0.825 ;
        RECT 1.010 0.645 2.220 0.695 ;
        RECT 0.515 0.305 1.775 0.475 ;
        RECT 1.945 0.280 2.220 0.645 ;
        RECT 2.455 0.085 2.625 0.525 ;
        RECT 2.795 0.280 3.135 0.695 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__o221ai_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o221ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.430 1.445 4.815 1.615 ;
        RECT 3.430 1.075 3.760 1.445 ;
        RECT 4.645 1.275 4.815 1.445 ;
        RECT 4.645 1.075 5.435 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.980 1.075 4.475 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.020 1.445 3.260 1.615 ;
        RECT 1.020 1.075 2.035 1.445 ;
        RECT 2.930 1.075 3.260 1.445 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.205 1.075 2.760 1.275 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.435 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.010 0.105 5.320 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.985500 ;
    PORT
      LAYER li1 ;
        RECT 0.560 1.955 0.810 2.465 ;
        RECT 2.340 1.955 2.590 2.125 ;
        RECT 4.100 1.955 4.350 2.125 ;
        RECT 0.560 1.785 4.350 1.955 ;
        RECT 0.560 1.445 0.850 1.785 ;
        RECT 0.605 0.865 0.850 1.445 ;
        RECT 0.520 0.645 0.850 0.865 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.140 1.455 0.390 2.635 ;
        RECT 0.980 2.125 1.750 2.635 ;
        RECT 1.920 2.295 3.010 2.465 ;
        RECT 1.920 2.125 2.170 2.295 ;
        RECT 2.760 2.125 3.010 2.295 ;
        RECT 3.180 2.125 3.510 2.635 ;
        RECT 3.680 2.295 4.770 2.465 ;
        RECT 3.680 2.125 3.930 2.295 ;
        RECT 4.520 1.785 4.770 2.295 ;
        RECT 4.985 1.455 5.190 2.635 ;
        RECT 0.100 0.475 0.350 0.895 ;
        RECT 1.020 0.645 3.050 0.905 ;
        RECT 3.220 0.735 5.230 0.905 ;
        RECT 1.020 0.475 1.270 0.645 ;
        RECT 3.220 0.475 3.550 0.735 ;
        RECT 4.060 0.725 5.230 0.735 ;
        RECT 0.100 0.255 1.270 0.475 ;
        RECT 1.460 0.255 3.550 0.475 ;
        RECT 3.720 0.085 3.890 0.555 ;
        RECT 4.060 0.255 4.390 0.725 ;
        RECT 4.560 0.085 4.730 0.555 ;
        RECT 4.900 0.255 5.230 0.725 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__o221ai_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o221ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o221ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 5.965 1.445 8.420 1.615 ;
        RECT 5.965 1.075 6.295 1.445 ;
        RECT 8.155 1.275 8.420 1.445 ;
        RECT 8.155 1.075 9.575 1.275 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.475 1.075 7.885 1.275 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 4.335 1.495 5.795 1.665 ;
        RECT 4.335 1.275 4.505 1.495 ;
        RECT 2.360 1.075 4.505 1.275 ;
        RECT 5.465 1.075 5.795 1.495 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 4.675 0.995 5.285 1.325 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 1.750 1.275 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.535 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.971000 ;
    PORT
      LAYER li1 ;
        RECT 0.575 1.615 0.825 2.465 ;
        RECT 1.415 1.955 1.665 2.465 ;
        RECT 3.995 2.005 4.285 2.125 ;
        RECT 4.875 2.005 5.085 2.125 ;
        RECT 6.675 2.005 6.885 2.125 ;
        RECT 3.995 1.955 6.885 2.005 ;
        RECT 7.475 1.955 7.725 2.125 ;
        RECT 1.415 1.615 2.125 1.955 ;
        RECT 3.995 1.835 7.725 1.955 ;
        RECT 3.995 1.615 4.165 1.835 ;
        RECT 5.965 1.785 7.725 1.835 ;
        RECT 0.575 1.445 4.165 1.615 ;
        RECT 1.920 0.865 2.125 1.445 ;
        RECT 0.535 0.645 2.125 0.865 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.155 1.485 0.405 2.635 ;
        RECT 0.995 1.825 1.245 2.635 ;
        RECT 1.835 2.125 2.605 2.635 ;
        RECT 2.775 1.955 3.025 2.465 ;
        RECT 3.195 2.125 3.445 2.635 ;
        RECT 3.615 2.295 5.585 2.465 ;
        RECT 3.615 1.955 3.825 2.295 ;
        RECT 4.455 2.175 4.705 2.295 ;
        RECT 5.255 2.175 5.585 2.295 ;
        RECT 5.755 2.175 6.005 2.635 ;
        RECT 6.175 2.295 8.145 2.465 ;
        RECT 6.175 2.175 6.505 2.295 ;
        RECT 7.055 2.125 7.305 2.295 ;
        RECT 2.775 1.785 3.825 1.955 ;
        RECT 7.895 1.955 8.145 2.295 ;
        RECT 8.315 2.125 8.565 2.635 ;
        RECT 8.735 1.955 8.985 2.465 ;
        RECT 7.895 1.785 8.985 1.955 ;
        RECT 8.735 1.445 8.985 1.785 ;
        RECT 9.155 1.445 9.405 2.635 ;
        RECT 0.115 0.475 0.365 0.895 ;
        RECT 5.465 0.820 9.445 0.905 ;
        RECT 2.315 0.735 9.445 0.820 ;
        RECT 2.315 0.645 6.085 0.735 ;
        RECT 0.115 0.255 5.585 0.475 ;
        RECT 5.755 0.255 6.085 0.645 ;
        RECT 6.595 0.725 7.765 0.735 ;
        RECT 6.255 0.085 6.425 0.555 ;
        RECT 6.595 0.255 6.925 0.725 ;
        RECT 7.095 0.085 7.265 0.555 ;
        RECT 7.435 0.255 7.765 0.725 ;
        RECT 8.275 0.725 9.445 0.735 ;
        RECT 7.935 0.085 8.105 0.555 ;
        RECT 8.275 0.255 8.605 0.725 ;
        RECT 8.775 0.085 8.945 0.555 ;
        RECT 9.115 0.255 9.445 0.725 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
  END
END sky130_fd_sc_hd__o221ai_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o311a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.995 1.280 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.520 1.325 1.790 2.070 ;
        RECT 1.450 0.995 1.790 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.980 1.325 2.215 2.070 ;
        RECT 1.980 0.995 2.270 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.440 0.995 2.840 1.325 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.350 0.995 3.595 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.105 3.675 1.015 ;
        RECT 0.140 -0.085 0.310 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.070 0.435 2.465 ;
        RECT 0.085 0.255 0.355 1.070 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.605 1.835 1.010 2.635 ;
        RECT 1.180 2.295 2.715 2.465 ;
        RECT 1.180 1.665 1.350 2.295 ;
        RECT 0.605 1.495 1.350 1.665 ;
        RECT 2.385 1.665 2.715 2.295 ;
        RECT 2.900 1.835 3.135 2.635 ;
        RECT 3.305 1.665 3.595 2.465 ;
        RECT 2.385 1.495 3.595 1.665 ;
        RECT 0.605 0.995 0.775 1.495 ;
        RECT 3.010 0.825 3.180 1.495 ;
        RECT 0.525 0.085 1.195 0.825 ;
        RECT 1.365 0.655 2.760 0.825 ;
        RECT 1.365 0.310 1.660 0.655 ;
        RECT 1.840 0.085 2.215 0.485 ;
        RECT 2.430 0.310 2.760 0.655 ;
        RECT 3.010 0.255 3.595 0.825 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__o311a_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o311a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.415 0.995 1.750 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.980 1.325 2.250 2.070 ;
        RECT 1.920 0.995 2.250 1.325 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.440 1.325 2.675 2.070 ;
        RECT 2.440 0.995 2.730 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.900 0.995 3.300 1.325 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.810 0.995 4.055 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.135 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.550 1.315 0.905 2.465 ;
        RECT 0.085 1.055 0.905 1.315 ;
        RECT 0.550 0.995 0.905 1.055 ;
        RECT 0.550 0.255 0.825 0.995 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 1.485 0.380 2.635 ;
        RECT 1.075 1.835 1.470 2.635 ;
        RECT 1.640 2.295 3.175 2.465 ;
        RECT 1.640 1.665 1.810 2.295 ;
        RECT 1.075 1.495 1.810 1.665 ;
        RECT 2.845 1.665 3.175 2.295 ;
        RECT 3.360 1.835 3.595 2.635 ;
        RECT 3.765 1.665 4.055 2.465 ;
        RECT 2.845 1.495 4.055 1.665 ;
        RECT 1.075 0.995 1.245 1.495 ;
        RECT 0.085 0.085 0.380 0.885 ;
        RECT 3.470 0.825 3.640 1.495 ;
        RECT 0.995 0.085 1.665 0.825 ;
        RECT 1.835 0.655 3.220 0.825 ;
        RECT 1.835 0.310 2.120 0.655 ;
        RECT 2.300 0.085 2.675 0.485 ;
        RECT 2.890 0.310 3.220 0.655 ;
        RECT 3.470 0.255 4.055 0.825 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__o311a_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o311a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.820 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 6.950 1.055 7.735 1.315 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 6.020 1.055 6.770 1.315 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.655 1.055 5.850 1.315 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.250 1.055 4.475 1.315 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.115 1.055 3.080 1.315 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.820 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.795 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.010 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.820 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.725 0.765 2.465 ;
        RECT 1.435 1.725 1.605 2.465 ;
        RECT 0.595 1.485 1.605 1.725 ;
        RECT 0.595 1.315 0.765 1.485 ;
        RECT 0.085 1.055 0.765 1.315 ;
        RECT 0.595 0.885 0.765 1.055 ;
        RECT 0.595 0.715 1.605 0.885 ;
        RECT 0.595 0.255 0.765 0.715 ;
        RECT 1.435 0.255 1.605 0.715 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.820 2.805 ;
        RECT 0.085 1.485 0.425 2.635 ;
        RECT 0.935 1.895 1.265 2.635 ;
        RECT 1.775 1.895 2.445 2.635 ;
        RECT 2.615 1.725 2.785 2.465 ;
        RECT 2.955 1.895 3.285 2.635 ;
        RECT 3.455 1.725 3.625 2.465 ;
        RECT 3.855 1.895 4.045 2.635 ;
        RECT 4.335 2.295 6.445 2.465 ;
        RECT 4.335 1.895 4.665 2.295 ;
        RECT 4.835 1.725 5.005 2.125 ;
        RECT 1.775 1.485 5.005 1.725 ;
        RECT 5.255 1.485 5.525 2.295 ;
        RECT 5.695 1.725 5.945 2.125 ;
        RECT 6.115 1.895 6.445 2.295 ;
        RECT 6.615 1.725 6.785 2.125 ;
        RECT 6.955 1.895 7.285 2.635 ;
        RECT 7.455 1.725 7.735 2.465 ;
        RECT 5.695 1.485 7.735 1.725 ;
        RECT 1.775 1.315 1.945 1.485 ;
        RECT 0.935 1.055 1.945 1.315 ;
        RECT 1.775 0.885 1.945 1.055 ;
        RECT 0.085 0.085 0.425 0.885 ;
        RECT 1.775 0.715 3.045 0.885 ;
        RECT 2.195 0.675 3.045 0.715 ;
        RECT 0.935 0.085 1.265 0.545 ;
        RECT 1.775 0.085 2.025 0.545 ;
        RECT 3.215 0.505 3.385 0.885 ;
        RECT 3.555 0.675 7.735 0.885 ;
        RECT 2.195 0.255 4.305 0.505 ;
        RECT 4.485 0.255 4.755 0.675 ;
        RECT 4.925 0.085 5.605 0.505 ;
        RECT 5.775 0.255 5.945 0.675 ;
        RECT 6.115 0.085 6.445 0.505 ;
        RECT 6.615 0.255 6.785 0.675 ;
        RECT 6.955 0.085 7.285 0.505 ;
        RECT 7.455 0.255 7.735 0.675 ;
        RECT 0.000 -0.085 7.820 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
  END
END sky130_fd_sc_hd__o311a_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o311ai_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.780 1.625 ;
        RECT 0.085 0.765 0.570 0.995 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.950 0.995 1.260 2.465 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.430 0.995 1.780 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.260 2.200 1.325 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.830 0.765 3.135 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.130 0.105 3.060 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.604000 ;
    PORT
      LAYER li1 ;
        RECT 1.430 1.665 1.980 2.465 ;
        RECT 2.650 1.665 3.135 2.465 ;
        RECT 1.430 1.495 3.135 1.665 ;
        RECT 2.445 0.595 2.660 1.495 ;
        RECT 2.445 0.255 3.135 0.595 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.795 0.780 2.635 ;
        RECT 2.150 1.835 2.480 2.635 ;
        RECT 0.740 0.655 1.750 0.825 ;
        RECT 0.085 0.085 0.570 0.595 ;
        RECT 0.740 0.255 0.910 0.655 ;
        RECT 1.080 0.085 1.410 0.485 ;
        RECT 1.580 0.255 1.750 0.655 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__o311ai_0

#--------EOF---------

MACRO sky130_fd_sc_hd__o311ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.780 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.950 0.995 1.260 2.465 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.430 0.995 1.780 1.325 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.985 0.320 2.200 1.325 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.830 0.995 3.135 1.325 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.130 0.105 3.060 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.942000 ;
    PORT
      LAYER li1 ;
        RECT 1.430 1.665 1.980 2.465 ;
        RECT 2.650 1.665 3.135 2.465 ;
        RECT 1.430 1.495 3.135 1.665 ;
        RECT 2.445 0.825 2.660 1.495 ;
        RECT 2.445 0.255 3.135 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.495 0.780 2.635 ;
        RECT 2.150 1.835 2.480 2.635 ;
        RECT 0.085 0.085 0.570 0.825 ;
        RECT 0.740 0.655 1.750 0.825 ;
        RECT 0.740 0.255 0.910 0.655 ;
        RECT 1.080 0.085 1.410 0.485 ;
        RECT 1.580 0.255 1.750 0.655 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__o311ai_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o311ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 1.105 1.315 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.275 1.055 2.155 1.315 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.325 1.055 3.075 1.315 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.365 1.055 4.385 1.315 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 5.085 1.055 5.895 1.315 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145 0.105 5.855 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.551000 ;
    PORT
      LAYER li1 ;
        RECT 2.415 1.725 2.665 2.125 ;
        RECT 3.335 1.725 3.505 2.465 ;
        RECT 4.515 1.725 4.825 2.465 ;
        RECT 5.495 1.725 5.895 2.465 ;
        RECT 2.415 1.485 5.895 1.725 ;
        RECT 4.555 0.885 4.915 1.485 ;
        RECT 4.555 0.655 5.895 0.885 ;
        RECT 5.515 0.255 5.895 0.655 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.085 1.725 0.465 2.465 ;
        RECT 0.635 1.895 0.965 2.635 ;
        RECT 1.135 1.725 1.305 2.465 ;
        RECT 1.475 2.295 3.165 2.465 ;
        RECT 1.475 1.895 1.805 2.295 ;
        RECT 1.975 1.725 2.225 2.125 ;
        RECT 2.835 1.895 3.165 2.295 ;
        RECT 3.675 1.895 4.345 2.635 ;
        RECT 4.995 1.895 5.325 2.635 ;
        RECT 0.085 1.485 2.225 1.725 ;
        RECT 0.085 0.655 4.385 0.885 ;
        RECT 0.085 0.255 0.485 0.655 ;
        RECT 0.655 0.085 0.985 0.485 ;
        RECT 1.155 0.255 1.325 0.655 ;
        RECT 1.495 0.085 1.825 0.485 ;
        RECT 1.995 0.255 2.165 0.655 ;
        RECT 2.335 0.085 3.105 0.485 ;
        RECT 3.275 0.255 3.445 0.655 ;
        RECT 3.615 0.255 5.345 0.485 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
  END
END sky130_fd_sc_hd__o311ai_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o311ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o311ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.055 1.775 1.315 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.945 1.055 3.615 1.315 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.805 1.055 5.885 1.315 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.055 1.055 7.695 1.315 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 7.865 1.055 9.090 1.315 ;
    END
  END C1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.065 0.105 9.595 1.015 ;
        RECT 0.125 -0.085 0.295 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.241000 ;
    PORT
      LAYER li1 ;
        RECT 4.055 1.725 4.305 2.115 ;
        RECT 4.975 1.725 5.145 2.115 ;
        RECT 5.815 1.725 6.005 2.465 ;
        RECT 6.675 1.725 6.845 2.465 ;
        RECT 7.515 1.725 7.685 2.465 ;
        RECT 8.355 1.725 8.525 2.465 ;
        RECT 9.195 1.725 9.575 2.465 ;
        RECT 4.055 1.485 9.575 1.725 ;
        RECT 9.260 0.885 9.575 1.485 ;
        RECT 7.895 0.655 9.575 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.085 1.725 0.405 2.465 ;
        RECT 0.595 1.895 0.925 2.635 ;
        RECT 1.095 1.725 1.265 2.465 ;
        RECT 1.435 1.895 1.765 2.635 ;
        RECT 1.935 1.725 2.105 2.465 ;
        RECT 2.275 2.295 5.645 2.465 ;
        RECT 2.275 1.895 2.605 2.295 ;
        RECT 2.775 1.725 2.945 2.115 ;
        RECT 3.115 1.895 3.445 2.295 ;
        RECT 3.615 1.725 3.865 2.115 ;
        RECT 4.475 1.895 4.805 2.295 ;
        RECT 5.315 1.895 5.645 2.295 ;
        RECT 6.175 1.895 6.505 2.635 ;
        RECT 7.015 1.895 7.345 2.635 ;
        RECT 7.855 1.895 8.185 2.635 ;
        RECT 8.695 1.895 9.025 2.635 ;
        RECT 0.085 1.485 3.865 1.725 ;
        RECT 0.085 0.085 0.505 0.885 ;
        RECT 0.675 0.655 7.385 0.885 ;
        RECT 0.675 0.255 0.845 0.655 ;
        RECT 1.015 0.085 1.345 0.485 ;
        RECT 1.515 0.255 1.685 0.655 ;
        RECT 1.855 0.085 2.185 0.485 ;
        RECT 2.355 0.255 2.525 0.655 ;
        RECT 2.695 0.085 3.025 0.485 ;
        RECT 3.195 0.255 3.365 0.655 ;
        RECT 3.535 0.085 3.885 0.485 ;
        RECT 4.055 0.255 4.225 0.655 ;
        RECT 4.395 0.085 4.725 0.485 ;
        RECT 4.895 0.255 5.065 0.655 ;
        RECT 7.555 0.485 7.725 0.885 ;
        RECT 5.235 0.085 5.585 0.485 ;
        RECT 5.755 0.255 9.575 0.485 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
  END
END sky130_fd_sc_hd__o311ai_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o2111a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111a_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.705 1.075 4.035 1.660 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.350 1.325 3.535 2.415 ;
        RECT 3.050 1.075 3.535 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.445 0.995 2.705 1.325 ;
        RECT 2.445 0.390 2.690 0.995 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.925 0.390 2.195 1.325 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.265 1.075 1.745 1.325 ;
        RECT 1.535 0.390 1.745 1.075 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.135 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.255 0.355 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.525 1.835 1.335 2.635 ;
        RECT 1.505 1.665 1.835 2.465 ;
        RECT 2.020 1.835 2.760 2.635 ;
        RECT 2.930 1.665 3.180 2.465 ;
        RECT 3.730 1.835 4.055 2.635 ;
        RECT 0.695 1.495 3.180 1.665 ;
        RECT 0.695 1.325 0.865 1.495 ;
        RECT 0.525 0.995 0.865 1.325 ;
        RECT 0.695 0.905 0.865 0.995 ;
        RECT 0.695 0.735 1.365 0.905 ;
        RECT 0.535 0.085 0.845 0.565 ;
        RECT 1.025 0.255 1.365 0.735 ;
        RECT 2.870 0.705 4.055 0.875 ;
        RECT 2.870 0.255 3.160 0.705 ;
        RECT 3.330 0.085 3.620 0.535 ;
        RECT 3.790 0.255 4.055 0.705 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__o2111a_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o2111a_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111a_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 4.310 1.315 4.515 2.355 ;
        RECT 3.830 1.005 4.515 1.315 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.370 1.325 3.660 2.370 ;
        RECT 3.300 0.995 3.660 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.680 1.075 3.100 1.615 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.005 0.255 2.390 1.615 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.075 1.835 1.615 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.305 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER li1 ;
        RECT 0.515 0.255 0.855 2.465 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.135 1.495 0.345 2.635 ;
        RECT 1.035 2.195 1.655 2.635 ;
        RECT 1.860 2.025 2.140 2.465 ;
        RECT 2.325 2.255 2.655 2.635 ;
        RECT 2.865 2.025 3.195 2.465 ;
        RECT 1.030 1.785 3.195 2.025 ;
        RECT 1.030 0.885 1.305 1.785 ;
        RECT 3.885 1.495 4.140 2.635 ;
        RECT 0.135 0.085 0.345 0.885 ;
        RECT 1.030 0.715 1.805 0.885 ;
        RECT 1.035 0.085 1.285 0.545 ;
        RECT 1.475 0.255 1.805 0.715 ;
        RECT 2.865 0.625 4.215 0.825 ;
        RECT 2.865 0.255 3.195 0.625 ;
        RECT 3.385 0.085 3.715 0.455 ;
        RECT 3.885 0.255 4.215 0.625 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__o2111a_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o2111a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111a_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.130 1.245 4.485 1.320 ;
        RECT 3.890 1.075 4.485 1.245 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.305 1.490 4.825 1.660 ;
        RECT 3.305 1.320 3.600 1.490 ;
        RECT 3.145 1.245 3.600 1.320 ;
        RECT 3.135 1.075 3.600 1.245 ;
        RECT 4.655 1.320 4.825 1.490 ;
        RECT 4.655 1.075 4.985 1.320 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.775 1.075 2.215 1.320 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.150 1.490 2.660 1.660 ;
        RECT 1.150 0.995 1.395 1.490 ;
        RECT 2.445 1.320 2.660 1.490 ;
        RECT 2.445 1.080 2.820 1.320 ;
        RECT 2.490 1.075 2.820 1.080 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.120 0.995 0.340 1.655 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 7.355 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.962500 ;
    PORT
      LAYER li1 ;
        RECT 5.755 1.665 5.925 2.465 ;
        RECT 6.585 1.665 6.775 2.465 ;
        RECT 5.755 1.495 7.275 1.665 ;
        RECT 7.005 0.865 7.275 1.495 ;
        RECT 5.650 0.695 7.275 0.865 ;
        RECT 5.650 0.255 5.875 0.695 ;
        RECT 6.545 0.255 6.745 0.695 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.090 2.005 0.345 2.465 ;
        RECT 0.515 2.175 0.845 2.635 ;
        RECT 1.015 2.005 1.230 2.465 ;
        RECT 1.400 2.175 1.625 2.635 ;
        RECT 1.795 2.005 2.025 2.465 ;
        RECT 2.195 2.175 2.525 2.635 ;
        RECT 2.695 2.005 3.285 2.465 ;
        RECT 3.805 2.180 4.135 2.635 ;
        RECT 4.775 2.005 5.065 2.465 ;
        RECT 5.245 2.170 5.585 2.635 ;
        RECT 0.090 2.000 5.065 2.005 ;
        RECT 0.090 1.835 5.550 2.000 ;
        RECT 6.095 1.835 6.415 2.635 ;
        RECT 6.945 1.835 7.270 2.635 ;
        RECT 0.515 1.830 5.550 1.835 ;
        RECT 0.100 0.485 0.345 0.825 ;
        RECT 0.515 0.655 0.860 1.830 ;
        RECT 5.380 1.320 5.550 1.830 ;
        RECT 5.380 1.075 6.760 1.320 ;
        RECT 1.720 0.655 4.795 0.885 ;
        RECT 0.100 0.255 2.940 0.485 ;
        RECT 3.110 0.085 3.440 0.485 ;
        RECT 3.610 0.255 3.825 0.655 ;
        RECT 3.995 0.085 4.365 0.485 ;
        RECT 4.535 0.255 4.795 0.655 ;
        RECT 5.035 0.085 5.300 0.545 ;
        RECT 6.075 0.085 6.375 0.525 ;
        RECT 6.915 0.085 7.275 0.525 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
  END
END sky130_fd_sc_hd__o2111a_4

#--------EOF---------

MACRO sky130_fd_sc_hd__o2111ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111ai_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.785 1.005 3.115 1.615 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.270 1.615 2.615 2.370 ;
        RECT 1.985 0.995 2.615 1.615 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.525 0.995 1.815 1.615 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.025 0.255 1.355 1.615 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.485 1.075 0.815 1.615 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.270 0.105 3.205 1.015 ;
        RECT 0.270 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.857250 ;
    PORT
      LAYER li1 ;
        RECT 0.790 2.025 1.025 2.465 ;
        RECT 1.750 2.025 2.095 2.465 ;
        RECT 0.085 1.785 2.095 2.025 ;
        RECT 0.085 0.885 0.315 1.785 ;
        RECT 0.085 0.255 0.690 0.885 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.290 2.195 0.620 2.635 ;
        RECT 1.210 2.255 1.540 2.635 ;
        RECT 2.785 1.795 3.115 2.635 ;
        RECT 1.750 0.625 3.115 0.825 ;
        RECT 1.750 0.255 2.095 0.625 ;
        RECT 2.285 0.085 2.615 0.455 ;
        RECT 2.785 0.255 3.115 0.625 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__o2111ai_1

#--------EOF---------

MACRO sky130_fd_sc_hd__o2111ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111ai_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 4.635 1.075 5.435 1.325 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 3.365 1.075 4.455 1.325 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 2.200 1.075 3.185 1.325 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 1.045 1.075 1.790 1.325 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.355 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.515 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.302000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.665 0.865 2.465 ;
        RECT 1.535 1.665 1.725 2.465 ;
        RECT 2.395 1.665 2.575 2.465 ;
        RECT 3.815 1.665 4.005 2.105 ;
        RECT 0.605 1.495 4.005 1.665 ;
        RECT 0.605 0.905 0.865 1.495 ;
        RECT 0.605 0.615 0.935 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.175 1.525 0.425 2.635 ;
        RECT 1.035 1.835 1.365 2.635 ;
        RECT 1.895 1.840 2.225 2.635 ;
        RECT 2.755 1.835 3.085 2.635 ;
        RECT 3.310 2.275 4.500 2.465 ;
        RECT 3.310 1.835 3.570 2.275 ;
        RECT 4.240 1.685 4.500 2.275 ;
        RECT 4.670 1.855 4.930 2.635 ;
        RECT 5.100 1.685 5.360 2.465 ;
        RECT 4.240 1.515 5.360 1.685 ;
        RECT 0.175 0.445 0.435 0.865 ;
        RECT 1.115 0.735 2.275 0.905 ;
        RECT 1.115 0.445 1.300 0.735 ;
        RECT 1.925 0.620 2.275 0.735 ;
        RECT 2.450 0.655 5.435 0.840 ;
        RECT 0.175 0.260 1.300 0.445 ;
        RECT 1.470 0.530 1.760 0.565 ;
        RECT 1.470 0.445 1.775 0.530 ;
        RECT 2.880 0.445 3.210 0.485 ;
        RECT 1.470 0.255 3.210 0.445 ;
        RECT 3.380 0.365 3.570 0.655 ;
        RECT 4.240 0.650 5.435 0.655 ;
        RECT 3.740 0.085 4.070 0.485 ;
        RECT 4.240 0.365 4.430 0.650 ;
        RECT 4.600 0.085 4.930 0.480 ;
        RECT 5.100 0.365 5.435 0.650 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__o2111ai_2

#--------EOF---------

MACRO sky130_fd_sc_hd__o2111ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__o2111ai_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 7.820 1.075 9.575 1.340 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 6.110 1.075 7.325 1.345 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 3.815 1.075 5.455 1.345 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.940 1.075 3.550 1.345 ;
    END
  END C1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.075 1.755 1.345 ;
    END
  END D1
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.530 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.984350 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.685 0.360 2.465 ;
        RECT 1.015 1.685 1.195 2.465 ;
        RECT 1.845 1.685 2.035 2.465 ;
        RECT 2.685 1.685 2.875 2.465 ;
        RECT 3.525 1.685 3.715 2.465 ;
        RECT 4.570 1.685 4.760 2.465 ;
        RECT 5.410 1.685 5.600 2.465 ;
        RECT 6.285 1.685 6.480 2.100 ;
        RECT 7.045 1.685 7.390 1.720 ;
        RECT 0.085 1.515 7.390 1.685 ;
        RECT 0.085 0.815 0.375 1.515 ;
        RECT 0.085 0.645 1.685 0.815 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.530 1.855 0.845 2.635 ;
        RECT 1.390 1.855 1.675 2.635 ;
        RECT 2.205 1.855 2.515 2.635 ;
        RECT 3.045 1.855 3.355 2.635 ;
        RECT 4.075 1.855 4.400 2.635 ;
        RECT 4.930 1.855 5.220 2.635 ;
        RECT 5.785 2.270 7.005 2.465 ;
        RECT 5.785 1.855 6.115 2.270 ;
        RECT 6.705 2.060 7.005 2.270 ;
        RECT 7.555 2.230 7.885 2.635 ;
        RECT 8.055 2.060 8.235 2.465 ;
        RECT 6.705 1.890 8.235 2.060 ;
        RECT 8.045 1.685 8.235 1.890 ;
        RECT 8.410 1.855 8.720 2.635 ;
        RECT 8.890 1.685 9.080 2.465 ;
        RECT 8.045 1.515 9.080 1.685 ;
        RECT 9.265 1.535 9.575 2.635 ;
        RECT 1.855 0.615 3.785 0.825 ;
        RECT 3.975 0.655 9.440 0.905 ;
        RECT 1.855 0.475 2.025 0.615 ;
        RECT 0.095 0.285 2.025 0.475 ;
        RECT 2.195 0.255 5.565 0.445 ;
        RECT 6.100 0.085 6.430 0.485 ;
        RECT 6.960 0.085 7.290 0.485 ;
        RECT 7.825 0.085 8.155 0.485 ;
        RECT 8.665 0.085 8.995 0.485 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
  END
END sky130_fd_sc_hd__o2111ai_4

#--------EOF---------

MACRO sky130_fd_sc_hd__or2_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.010 0.995 1.335 1.615 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.995 0.500 1.615 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150 0.335 1.985 1.015 ;
        RECT 0.150 0.085 0.315 0.335 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.326800 ;
    PORT
      LAYER li1 ;
        RECT 1.645 2.135 2.180 2.465 ;
        RECT 1.865 0.825 2.180 2.135 ;
        RECT 1.565 0.525 2.180 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.270 1.955 0.660 2.130 ;
        RECT 1.145 2.125 1.475 2.635 ;
        RECT 0.270 1.785 1.695 1.955 ;
        RECT 0.670 0.825 0.840 1.785 ;
        RECT 1.525 0.995 1.695 1.785 ;
        RECT 0.250 0.085 0.490 0.825 ;
        RECT 0.670 0.425 0.950 0.825 ;
        RECT 1.180 0.085 1.395 0.825 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__or2_0

#--------EOF---------

MACRO sky130_fd_sc_hd__or2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.010 0.765 1.275 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.765 0.500 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.055 0.785 1.985 1.015 ;
        RECT 0.150 0.105 1.985 0.785 ;
        RECT 0.150 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.509000 ;
    PORT
      LAYER li1 ;
        RECT 1.645 1.845 2.180 2.465 ;
        RECT 1.865 0.825 2.180 1.845 ;
        RECT 1.565 0.255 2.180 0.825 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.270 1.665 0.660 1.840 ;
        RECT 1.145 1.835 1.475 2.635 ;
        RECT 0.270 1.495 1.695 1.665 ;
        RECT 0.670 0.595 0.840 1.495 ;
        RECT 1.525 0.995 1.695 1.495 ;
        RECT 0.250 0.085 0.490 0.595 ;
        RECT 0.670 0.265 0.950 0.595 ;
        RECT 1.180 0.085 1.395 0.595 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__or2_1

#--------EOF---------

MACRO sky130_fd_sc_hd__or2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.865 0.765 1.275 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.150 0.765 0.345 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.910 0.785 2.280 1.015 ;
        RECT 0.005 0.105 2.280 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 1.440 2.005 1.770 2.465 ;
        RECT 1.440 1.835 2.215 2.005 ;
        RECT 1.785 0.825 2.215 1.835 ;
        RECT 1.520 0.655 2.215 0.825 ;
        RECT 1.520 0.385 1.690 0.655 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.155 1.665 0.515 1.840 ;
        RECT 1.100 1.835 1.270 2.635 ;
        RECT 1.940 2.175 2.110 2.635 ;
        RECT 0.155 1.495 1.615 1.665 ;
        RECT 0.515 0.595 0.695 1.495 ;
        RECT 1.445 0.995 1.615 1.495 ;
        RECT 0.105 0.085 0.345 0.595 ;
        RECT 0.515 0.255 0.805 0.595 ;
        RECT 1.035 0.085 1.350 0.595 ;
        RECT 1.860 0.085 2.190 0.485 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__or2_2

#--------EOF---------

MACRO sky130_fd_sc_hd__or2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.865 0.995 1.240 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.765 0.345 1.325 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 3.120 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 1.440 2.005 1.770 2.465 ;
        RECT 2.280 2.005 2.610 2.465 ;
        RECT 1.440 1.835 2.610 2.005 ;
        RECT 2.280 1.665 2.610 1.835 ;
        RECT 2.280 1.495 3.135 1.665 ;
        RECT 2.790 0.905 3.135 1.495 ;
        RECT 1.440 0.735 3.135 0.905 ;
        RECT 1.440 0.265 1.770 0.735 ;
        RECT 2.280 0.265 2.610 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.155 1.665 0.515 2.465 ;
        RECT 1.060 1.835 1.230 2.635 ;
        RECT 1.940 2.175 2.110 2.635 ;
        RECT 2.780 1.835 2.950 2.635 ;
        RECT 0.155 1.495 1.615 1.665 ;
        RECT 0.515 0.825 0.695 1.495 ;
        RECT 1.410 1.245 1.615 1.495 ;
        RECT 1.410 1.075 2.620 1.245 ;
        RECT 0.105 0.085 0.345 0.595 ;
        RECT 0.515 0.290 0.845 0.825 ;
        RECT 1.060 0.085 1.230 0.825 ;
        RECT 1.940 0.085 2.110 0.565 ;
        RECT 2.780 0.085 2.950 0.565 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__or2_4

#--------EOF---------

MACRO sky130_fd_sc_hd__or2b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.540 2.085 1.735 2.415 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.425 1.325 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.810 0.815 2.755 1.015 ;
        RECT 0.005 0.135 2.755 0.815 ;
        RECT 0.150 -0.085 0.320 0.135 ;
        RECT 1.810 0.105 2.755 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.495 2.675 2.465 ;
        RECT 2.505 0.760 2.675 1.495 ;
        RECT 2.405 0.415 2.675 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.090 1.495 0.345 2.635 ;
        RECT 0.595 1.325 0.765 1.885 ;
        RECT 0.990 1.665 1.410 1.915 ;
        RECT 1.915 1.835 2.195 2.635 ;
        RECT 0.990 1.495 2.235 1.665 ;
        RECT 2.065 1.325 2.235 1.495 ;
        RECT 0.595 0.995 1.335 1.325 ;
        RECT 2.065 0.995 2.295 1.325 ;
        RECT 0.595 0.905 0.845 0.995 ;
        RECT 0.110 0.735 0.845 0.905 ;
        RECT 2.065 0.825 2.235 0.995 ;
        RECT 0.110 0.265 0.420 0.735 ;
        RECT 1.495 0.655 2.235 0.825 ;
        RECT 0.590 0.085 1.325 0.565 ;
        RECT 1.495 0.305 1.665 0.655 ;
        RECT 1.835 0.085 2.215 0.485 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__or2b_1

#--------EOF---------

MACRO sky130_fd_sc_hd__or2b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.540 2.085 1.730 2.415 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.325 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.805 0.815 3.210 1.015 ;
        RECT 0.005 0.135 3.210 0.815 ;
        RECT 0.145 -0.085 0.315 0.135 ;
        RECT 1.805 0.105 3.210 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 2.400 1.495 2.630 2.465 ;
        RECT 2.460 0.760 2.630 1.495 ;
        RECT 2.400 0.415 2.630 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 0.595 1.325 0.765 1.885 ;
        RECT 0.985 1.665 1.405 1.915 ;
        RECT 1.910 1.835 2.190 2.635 ;
        RECT 0.985 1.495 2.230 1.665 ;
        RECT 2.060 1.325 2.230 1.495 ;
        RECT 2.800 1.460 3.055 2.635 ;
        RECT 0.595 0.995 1.330 1.325 ;
        RECT 2.060 0.995 2.290 1.325 ;
        RECT 0.595 0.905 0.840 0.995 ;
        RECT 0.105 0.735 0.840 0.905 ;
        RECT 2.060 0.825 2.230 0.995 ;
        RECT 0.105 0.265 0.420 0.735 ;
        RECT 1.490 0.655 2.230 0.825 ;
        RECT 0.590 0.085 1.320 0.565 ;
        RECT 1.490 0.305 1.660 0.655 ;
        RECT 1.830 0.085 2.210 0.485 ;
        RECT 2.800 0.085 3.055 0.925 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__or2b_2

#--------EOF---------

MACRO sky130_fd_sc_hd__or2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or2b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.630 1.075 2.320 1.275 ;
    END
  END A
  PIN B_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.425 1.955 ;
    END
  END B_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.780 0.815 4.075 1.015 ;
        RECT 0.005 0.135 4.075 0.815 ;
        RECT 0.145 0.105 4.075 0.135 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 2.365 1.955 2.615 2.465 ;
        RECT 3.205 1.955 3.455 2.465 ;
        RECT 2.365 1.785 3.455 1.955 ;
        RECT 2.830 1.615 3.455 1.785 ;
        RECT 2.830 1.445 4.055 1.615 ;
        RECT 3.670 0.905 4.055 1.445 ;
        RECT 2.325 0.735 4.055 0.905 ;
        RECT 2.325 0.290 2.655 0.735 ;
        RECT 3.165 0.290 3.495 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.090 2.125 0.345 2.635 ;
        RECT 0.595 1.325 0.765 2.465 ;
        RECT 0.990 1.615 1.460 2.465 ;
        RECT 1.915 1.835 2.195 2.635 ;
        RECT 2.785 2.135 3.035 2.635 ;
        RECT 3.625 1.795 3.875 2.635 ;
        RECT 0.990 1.495 2.660 1.615 ;
        RECT 1.290 1.445 2.660 1.495 ;
        RECT 0.595 0.995 1.120 1.325 ;
        RECT 0.595 0.905 0.845 0.995 ;
        RECT 0.110 0.735 0.845 0.905 ;
        RECT 1.290 0.905 1.460 1.445 ;
        RECT 2.490 1.245 2.660 1.445 ;
        RECT 2.490 1.075 3.500 1.245 ;
        RECT 1.290 0.735 1.745 0.905 ;
        RECT 0.110 0.265 0.420 0.735 ;
        RECT 0.590 0.085 1.245 0.565 ;
        RECT 1.415 0.305 1.745 0.735 ;
        RECT 1.980 0.085 2.155 0.905 ;
        RECT 2.825 0.085 2.995 0.550 ;
        RECT 3.665 0.085 3.835 0.550 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__or2b_4

#--------EOF---------

MACRO sky130_fd_sc_hd__or3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.300 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.600 1.325 0.795 1.615 ;
        RECT 0.600 0.995 1.425 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.125 1.275 2.415 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.430 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.300 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.340 0.815 2.295 1.015 ;
        RECT 0.015 0.135 2.295 0.815 ;
        RECT 0.140 -0.085 0.310 0.135 ;
        RECT 1.340 0.105 2.295 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.490 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.300 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER li1 ;
        RECT 1.935 1.495 2.210 2.465 ;
        RECT 2.040 0.760 2.210 1.495 ;
        RECT 1.935 0.415 2.210 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.300 2.805 ;
        RECT 0.105 1.785 1.275 1.955 ;
        RECT 1.445 1.835 1.725 2.635 ;
        RECT 0.105 1.495 0.430 1.785 ;
        RECT 1.105 1.665 1.275 1.785 ;
        RECT 1.105 1.495 1.765 1.665 ;
        RECT 1.595 1.325 1.765 1.495 ;
        RECT 1.595 0.995 1.870 1.325 ;
        RECT 1.595 0.825 1.765 0.995 ;
        RECT 0.100 0.655 1.765 0.825 ;
        RECT 0.100 0.305 0.355 0.655 ;
        RECT 0.525 0.085 0.855 0.485 ;
        RECT 1.025 0.305 1.195 0.655 ;
        RECT 1.365 0.085 1.745 0.485 ;
        RECT 0.000 -0.085 2.300 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
  END
END sky130_fd_sc_hd__or3_1

#--------EOF---------

MACRO sky130_fd_sc_hd__or3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.605 1.325 0.830 1.615 ;
        RECT 0.605 0.995 1.430 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.125 1.280 2.415 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.995 0.435 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.345 0.815 2.725 1.015 ;
        RECT 0.020 0.135 2.725 0.815 ;
        RECT 0.145 -0.085 0.315 0.135 ;
        RECT 1.345 0.105 2.725 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 1.940 1.495 2.215 2.465 ;
        RECT 2.045 0.760 2.215 1.495 ;
        RECT 1.940 0.415 2.215 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.105 1.785 1.270 1.955 ;
        RECT 1.450 1.835 1.730 2.635 ;
        RECT 0.105 1.495 0.435 1.785 ;
        RECT 1.100 1.665 1.270 1.785 ;
        RECT 1.100 1.495 1.770 1.665 ;
        RECT 1.600 1.325 1.770 1.495 ;
        RECT 2.385 1.430 2.675 2.635 ;
        RECT 1.600 0.995 1.875 1.325 ;
        RECT 1.600 0.825 1.770 0.995 ;
        RECT 0.105 0.655 1.770 0.825 ;
        RECT 0.105 0.305 0.360 0.655 ;
        RECT 0.530 0.085 0.860 0.485 ;
        RECT 1.030 0.305 1.200 0.655 ;
        RECT 1.370 0.085 1.750 0.485 ;
        RECT 2.385 0.085 2.675 0.915 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__or3_2

#--------EOF---------

MACRO sky130_fd_sc_hd__or3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.225 1.075 1.700 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.595 1.325 0.830 2.050 ;
        RECT 0.595 1.075 1.055 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.040 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 2.345 1.625 2.595 2.465 ;
        RECT 3.185 1.625 3.435 2.465 ;
        RECT 2.345 1.455 4.055 1.625 ;
        RECT 3.765 0.905 4.055 1.455 ;
        RECT 2.305 0.735 4.055 0.905 ;
        RECT 2.305 0.265 2.635 0.735 ;
        RECT 3.145 0.265 3.475 0.735 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 2.295 1.265 2.465 ;
        RECT 0.085 1.495 0.425 2.295 ;
        RECT 1.000 1.665 1.265 2.295 ;
        RECT 1.435 1.835 2.135 2.635 ;
        RECT 2.765 1.795 3.015 2.635 ;
        RECT 3.605 1.795 3.855 2.635 ;
        RECT 1.000 1.495 2.090 1.665 ;
        RECT 1.870 1.245 2.090 1.495 ;
        RECT 1.870 1.075 3.595 1.245 ;
        RECT 1.870 0.905 2.090 1.075 ;
        RECT 0.085 0.725 2.090 0.905 ;
        RECT 0.085 0.255 0.425 0.725 ;
        RECT 0.595 0.085 0.765 0.555 ;
        RECT 0.935 0.255 1.265 0.725 ;
        RECT 1.435 0.085 2.135 0.555 ;
        RECT 2.805 0.085 2.975 0.555 ;
        RECT 3.645 0.085 3.815 0.555 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__or3_4

#--------EOF---------

MACRO sky130_fd_sc_hd__or3b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.525 1.325 1.770 1.615 ;
        RECT 1.525 0.995 2.350 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.585 2.125 2.200 2.455 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 1.075 0.425 1.325 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.815 0.935 1.015 ;
        RECT 2.270 0.815 3.215 1.015 ;
        RECT 0.005 0.335 3.215 0.815 ;
        RECT 0.145 0.135 3.215 0.335 ;
        RECT 0.145 -0.085 0.315 0.135 ;
        RECT 2.270 0.105 3.215 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.453750 ;
    PORT
      LAYER li1 ;
        RECT 2.860 1.495 3.135 2.465 ;
        RECT 2.965 0.760 3.135 1.495 ;
        RECT 2.860 0.415 3.135 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.495 0.345 2.635 ;
        RECT 0.595 1.325 0.765 1.885 ;
        RECT 1.025 1.785 2.200 1.955 ;
        RECT 2.370 1.835 2.650 2.635 ;
        RECT 1.025 1.495 1.355 1.785 ;
        RECT 2.030 1.665 2.200 1.785 ;
        RECT 2.030 1.495 2.690 1.665 ;
        RECT 2.520 1.325 2.690 1.495 ;
        RECT 0.595 0.995 1.310 1.325 ;
        RECT 2.520 0.995 2.795 1.325 ;
        RECT 0.595 0.905 0.845 0.995 ;
        RECT 0.085 0.085 0.345 0.905 ;
        RECT 0.515 0.485 0.845 0.905 ;
        RECT 2.520 0.825 2.690 0.995 ;
        RECT 1.025 0.655 2.690 0.825 ;
        RECT 1.025 0.255 1.285 0.655 ;
        RECT 1.455 0.085 1.785 0.485 ;
        RECT 1.955 0.305 2.125 0.655 ;
        RECT 2.295 0.085 2.670 0.485 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__or3b_1

#--------EOF---------

MACRO sky130_fd_sc_hd__or3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.695 1.075 2.230 1.615 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.935 2.125 3.135 2.365 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.640 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.490 0.815 1.845 1.015 ;
        RECT 0.490 0.785 3.170 0.815 ;
        RECT 0.005 0.135 3.170 0.785 ;
        RECT 0.005 0.105 1.845 0.135 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.935 1.495 1.330 1.700 ;
        RECT 0.935 0.595 1.105 1.495 ;
        RECT 0.935 0.265 1.285 0.595 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 2.040 0.345 2.220 ;
        RECT 0.550 2.210 0.910 2.635 ;
        RECT 1.425 2.210 1.755 2.635 ;
        RECT 0.085 1.955 1.720 2.040 ;
        RECT 0.085 1.870 2.660 1.955 ;
        RECT 0.085 1.810 0.765 1.870 ;
        RECT 0.595 0.905 0.765 1.810 ;
        RECT 1.550 1.785 2.660 1.870 ;
        RECT 2.490 1.325 2.660 1.785 ;
        RECT 2.830 1.495 3.135 1.925 ;
        RECT 0.085 0.735 0.765 0.905 ;
        RECT 1.275 0.935 1.445 1.325 ;
        RECT 2.490 0.995 2.790 1.325 ;
        RECT 1.275 0.905 1.595 0.935 ;
        RECT 1.275 0.825 2.160 0.905 ;
        RECT 2.965 0.825 3.135 1.495 ;
        RECT 1.275 0.765 3.135 0.825 ;
        RECT 1.425 0.735 3.135 0.765 ;
        RECT 0.085 0.290 0.345 0.735 ;
        RECT 1.990 0.655 3.135 0.735 ;
        RECT 0.595 0.085 0.765 0.565 ;
        RECT 1.520 0.085 1.690 0.565 ;
        RECT 1.990 0.305 2.160 0.655 ;
        RECT 2.830 0.605 3.135 0.655 ;
        RECT 2.330 0.085 2.660 0.485 ;
        RECT 2.830 0.305 3.085 0.605 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__or3b_2

#--------EOF---------

MACRO sky130_fd_sc_hd__or3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or3b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.400 1.415 2.720 1.700 ;
        RECT 2.535 0.995 2.720 1.415 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.890 0.995 3.200 1.700 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.640 ;
    END
  END C_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.490 0.785 4.000 1.015 ;
        RECT 0.005 0.105 4.000 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.935 1.415 2.220 1.700 ;
        RECT 0.935 0.905 1.105 1.415 ;
        RECT 0.935 0.735 2.025 0.905 ;
        RECT 1.000 0.285 1.330 0.735 ;
        RECT 1.855 0.585 2.025 0.735 ;
        RECT 1.855 0.255 2.090 0.585 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 2.040 0.345 2.220 ;
        RECT 0.550 2.210 0.910 2.635 ;
        RECT 1.420 2.210 1.750 2.635 ;
        RECT 2.255 2.210 2.595 2.635 ;
        RECT 3.520 2.210 4.055 2.425 ;
        RECT 0.085 1.870 3.620 2.040 ;
        RECT 0.085 1.810 0.765 1.870 ;
        RECT 0.595 0.905 0.765 1.810 ;
        RECT 3.390 1.325 3.620 1.870 ;
        RECT 1.275 1.075 2.365 1.245 ;
        RECT 0.085 0.735 0.765 0.905 ;
        RECT 2.195 0.890 2.365 1.075 ;
        RECT 3.390 0.995 3.680 1.325 ;
        RECT 2.195 0.825 2.400 0.890 ;
        RECT 3.850 0.825 4.055 2.210 ;
        RECT 0.085 0.290 0.345 0.735 ;
        RECT 2.195 0.720 4.055 0.825 ;
        RECT 2.250 0.655 4.055 0.720 ;
        RECT 0.620 0.085 0.790 0.565 ;
        RECT 1.500 0.085 1.670 0.565 ;
        RECT 2.260 0.085 2.590 0.485 ;
        RECT 2.760 0.305 2.930 0.655 ;
        RECT 3.660 0.605 4.055 0.655 ;
        RECT 3.100 0.085 3.490 0.485 ;
        RECT 3.660 0.305 3.915 0.605 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__or3b_4

#--------EOF---------

MACRO sky130_fd_sc_hd__or4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.490 0.995 1.895 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 2.125 1.745 2.415 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.610 0.995 1.320 1.615 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.090 0.755 0.440 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.810 0.815 2.755 1.015 ;
        RECT 0.005 0.135 2.755 0.815 ;
        RECT 0.150 -0.085 0.320 0.135 ;
        RECT 1.810 0.105 2.755 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 2.950 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.495 2.675 2.465 ;
        RECT 2.505 0.760 2.675 1.495 ;
        RECT 2.405 0.415 2.675 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 2.760 2.805 ;
        RECT 0.090 1.785 1.680 1.955 ;
        RECT 1.915 1.835 2.195 2.635 ;
        RECT 0.090 1.495 0.410 1.785 ;
        RECT 1.510 1.665 1.680 1.785 ;
        RECT 1.510 1.495 2.235 1.665 ;
        RECT 2.065 1.325 2.235 1.495 ;
        RECT 2.065 0.995 2.335 1.325 ;
        RECT 2.065 0.825 2.235 0.995 ;
        RECT 0.625 0.655 2.235 0.825 ;
        RECT 0.095 0.085 0.425 0.585 ;
        RECT 0.625 0.305 0.795 0.655 ;
        RECT 0.995 0.085 1.325 0.485 ;
        RECT 1.495 0.305 1.665 0.655 ;
        RECT 1.835 0.085 2.215 0.485 ;
        RECT 0.000 -0.085 2.760 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
  END
END sky130_fd_sc_hd__or4_1

#--------EOF---------

MACRO sky130_fd_sc_hd__or4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.490 0.995 1.895 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 2.125 1.745 2.415 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.610 0.995 1.320 1.615 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.755 0.440 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 1.810 0.815 3.210 1.015 ;
        RECT 0.005 0.135 3.210 0.815 ;
        RECT 0.150 -0.085 0.320 0.135 ;
        RECT 1.810 0.105 3.210 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 2.405 1.495 2.680 2.465 ;
        RECT 2.510 0.760 2.680 1.495 ;
        RECT 2.405 0.415 2.680 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.785 1.680 1.955 ;
        RECT 1.915 1.835 2.195 2.635 ;
        RECT 0.085 1.495 0.410 1.785 ;
        RECT 1.510 1.665 1.680 1.785 ;
        RECT 1.510 1.495 2.235 1.665 ;
        RECT 2.065 1.325 2.235 1.495 ;
        RECT 2.850 1.455 3.020 2.635 ;
        RECT 2.065 0.995 2.340 1.325 ;
        RECT 2.065 0.825 2.235 0.995 ;
        RECT 0.625 0.655 2.235 0.825 ;
        RECT 0.090 0.085 0.425 0.585 ;
        RECT 0.625 0.305 0.795 0.655 ;
        RECT 0.995 0.085 1.325 0.485 ;
        RECT 1.495 0.305 1.665 0.655 ;
        RECT 1.835 0.085 2.215 0.485 ;
        RECT 2.850 0.085 3.020 1.000 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__or4_2

#--------EOF---------

MACRO sky130_fd_sc_hd__or4_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.840 1.445 2.275 1.615 ;
        RECT 1.840 0.995 2.010 1.445 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.400 1.785 1.720 2.375 ;
        RECT 1.400 1.450 1.610 1.785 ;
        RECT 1.280 0.995 1.610 1.450 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.880 1.620 1.230 2.375 ;
        RECT 0.880 0.995 1.050 1.620 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.755 0.370 1.325 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.030 0.105 4.135 1.015 ;
        RECT 0.140 -0.085 0.310 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 2.480 1.625 2.730 2.465 ;
        RECT 3.320 1.625 3.570 2.465 ;
        RECT 2.480 1.455 4.055 1.625 ;
        RECT 3.810 0.905 4.055 1.455 ;
        RECT 2.520 0.725 4.055 0.905 ;
        RECT 2.520 0.255 2.770 0.725 ;
        RECT 3.280 0.255 3.610 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.115 1.665 0.450 2.450 ;
        RECT 2.005 1.795 2.255 2.635 ;
        RECT 2.900 1.795 3.150 2.635 ;
        RECT 3.740 1.795 3.990 2.635 ;
        RECT 0.115 1.495 0.710 1.665 ;
        RECT 0.540 0.825 0.710 1.495 ;
        RECT 2.180 1.075 3.640 1.245 ;
        RECT 2.180 0.825 2.350 1.075 ;
        RECT 0.540 0.655 2.350 0.825 ;
        RECT 0.120 0.085 0.370 0.585 ;
        RECT 0.700 0.305 0.870 0.655 ;
        RECT 1.070 0.085 1.400 0.485 ;
        RECT 1.570 0.305 1.740 0.655 ;
        RECT 1.960 0.085 2.340 0.485 ;
        RECT 2.940 0.085 3.110 0.555 ;
        RECT 3.780 0.085 3.950 0.555 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__or4_4

#--------EOF---------

MACRO sky130_fd_sc_hd__or4b_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4b_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.430 0.995 2.810 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.610 2.125 2.660 2.415 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.520 0.995 2.260 1.615 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.755 0.425 1.325 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.725 0.815 3.675 1.015 ;
        RECT 0.005 0.135 3.675 0.815 ;
        RECT 0.150 -0.085 0.320 0.135 ;
        RECT 2.725 0.105 3.675 0.135 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.453750 ;
    PORT
      LAYER li1 ;
        RECT 3.320 1.495 3.595 2.465 ;
        RECT 3.425 0.760 3.595 1.495 ;
        RECT 3.320 0.415 3.595 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.085 1.560 0.425 2.635 ;
        RECT 0.595 1.325 0.835 1.920 ;
        RECT 1.030 1.785 2.660 1.955 ;
        RECT 2.830 1.835 3.110 2.635 ;
        RECT 1.030 1.495 1.350 1.785 ;
        RECT 2.490 1.665 2.660 1.785 ;
        RECT 2.490 1.495 3.150 1.665 ;
        RECT 2.980 1.325 3.150 1.495 ;
        RECT 0.595 0.995 1.250 1.325 ;
        RECT 2.980 0.995 3.255 1.325 ;
        RECT 0.085 0.085 0.425 0.585 ;
        RECT 0.595 0.305 0.840 0.995 ;
        RECT 2.980 0.825 3.150 0.995 ;
        RECT 1.565 0.655 3.150 0.825 ;
        RECT 1.035 0.085 1.365 0.585 ;
        RECT 1.565 0.305 1.735 0.655 ;
        RECT 1.910 0.085 2.240 0.485 ;
        RECT 2.410 0.305 2.580 0.655 ;
        RECT 2.750 0.085 3.130 0.485 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__or4b_1

#--------EOF---------

MACRO sky130_fd_sc_hd__or4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4b_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.755 1.075 2.320 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 1.985 2.125 2.670 2.415 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.550 1.075 3.550 1.275 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.075 0.425 1.435 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.490 0.815 1.840 1.015 ;
        RECT 0.005 0.135 3.645 0.815 ;
        RECT 0.150 0.105 1.840 0.135 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.870 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.935 1.495 1.250 1.825 ;
        RECT 0.935 0.790 1.105 1.495 ;
        RECT 0.935 0.680 1.245 0.790 ;
        RECT 0.935 0.675 1.250 0.680 ;
        RECT 0.970 0.260 1.250 0.675 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.680 2.805 ;
        RECT 0.515 2.335 0.845 2.635 ;
        RECT 1.480 2.335 1.815 2.635 ;
        RECT 2.860 2.215 3.345 2.385 ;
        RECT 0.510 1.995 1.715 2.165 ;
        RECT 0.510 1.890 0.765 1.995 ;
        RECT 0.085 1.605 0.765 1.890 ;
        RECT 1.440 1.955 1.715 1.995 ;
        RECT 2.860 1.955 3.030 2.215 ;
        RECT 1.440 1.785 3.030 1.955 ;
        RECT 3.225 1.615 3.560 1.815 ;
        RECT 0.595 0.905 0.765 1.605 ;
        RECT 1.420 1.450 3.560 1.615 ;
        RECT 1.415 1.445 3.560 1.450 ;
        RECT 1.415 1.425 1.665 1.445 ;
        RECT 1.415 1.420 1.655 1.425 ;
        RECT 1.415 1.410 1.645 1.420 ;
        RECT 1.415 1.400 1.630 1.410 ;
        RECT 1.415 1.390 1.625 1.400 ;
        RECT 1.415 1.380 1.620 1.390 ;
        RECT 1.415 1.370 1.610 1.380 ;
        RECT 1.415 1.355 1.600 1.370 ;
        RECT 1.415 1.325 1.585 1.355 ;
        RECT 1.290 0.995 1.585 1.325 ;
        RECT 0.085 0.735 0.765 0.905 ;
        RECT 1.415 0.905 1.585 0.995 ;
        RECT 1.415 0.735 3.055 0.905 ;
        RECT 0.085 0.325 0.350 0.735 ;
        RECT 0.630 0.085 0.800 0.565 ;
        RECT 1.435 0.085 1.815 0.485 ;
        RECT 1.985 0.305 2.155 0.735 ;
        RECT 2.385 0.085 2.715 0.485 ;
        RECT 2.885 0.305 3.055 0.735 ;
        RECT 3.225 0.085 3.555 0.585 ;
        RECT 0.000 -0.085 3.680 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
  END
END sky130_fd_sc_hd__or4b_2

#--------EOF---------

MACRO sky130_fd_sc_hd__or4b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4b_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.755 1.445 3.190 1.615 ;
        RECT 2.755 0.995 2.925 1.445 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.335 1.785 2.635 2.375 ;
        RECT 2.335 1.450 2.525 1.785 ;
        RECT 2.195 0.995 2.525 1.450 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 1.795 1.620 2.155 2.375 ;
        RECT 1.795 0.995 1.965 1.620 ;
    END
  END C
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.105 0.995 0.445 1.955 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.335 5.050 1.015 ;
        RECT 0.145 0.105 5.050 0.335 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 3.395 1.625 3.645 2.465 ;
        RECT 4.235 1.625 4.485 2.465 ;
        RECT 3.395 1.455 4.965 1.625 ;
        RECT 4.725 0.905 4.965 1.455 ;
        RECT 3.435 0.725 4.965 0.905 ;
        RECT 3.435 0.255 3.685 0.725 ;
        RECT 4.195 0.255 4.525 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 0.085 2.135 0.365 2.635 ;
        RECT 0.595 2.065 0.785 2.455 ;
        RECT 0.615 1.325 0.785 2.065 ;
        RECT 1.035 1.745 1.365 2.450 ;
        RECT 2.920 1.795 3.170 2.635 ;
        RECT 3.815 1.795 4.065 2.635 ;
        RECT 4.655 1.795 4.905 2.635 ;
        RECT 1.035 1.575 1.625 1.745 ;
        RECT 0.615 0.995 1.215 1.325 ;
        RECT 0.615 0.905 0.785 0.995 ;
        RECT 0.085 0.085 0.345 0.825 ;
        RECT 0.595 0.435 0.785 0.905 ;
        RECT 1.455 0.825 1.625 1.575 ;
        RECT 3.095 1.075 4.555 1.245 ;
        RECT 3.095 0.825 3.265 1.075 ;
        RECT 1.455 0.655 3.265 0.825 ;
        RECT 1.035 0.085 1.285 0.585 ;
        RECT 1.615 0.305 1.785 0.655 ;
        RECT 1.985 0.085 2.315 0.485 ;
        RECT 2.485 0.305 2.655 0.655 ;
        RECT 2.875 0.085 3.255 0.485 ;
        RECT 3.855 0.085 4.025 0.555 ;
        RECT 4.695 0.085 4.865 0.555 ;
        RECT 0.000 -0.085 5.060 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
  END
END sky130_fd_sc_hd__or4b_4

#--------EOF---------

MACRO sky130_fd_sc_hd__or4bb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4bb_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.615 0.995 3.270 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.480 2.125 3.120 2.455 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.695 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.995 1.235 1.325 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.040 0.785 1.415 1.015 ;
        RECT 3.185 0.785 4.135 1.015 ;
        RECT 0.040 0.335 4.135 0.785 ;
        RECT 0.145 -0.085 0.315 0.335 ;
        RECT 1.425 0.105 4.135 0.335 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.453750 ;
    PORT
      LAYER li1 ;
        RECT 3.780 1.495 4.055 2.465 ;
        RECT 3.885 0.760 4.055 1.495 ;
        RECT 3.780 0.415 4.055 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 2.035 0.345 2.455 ;
        RECT 0.515 2.205 0.845 2.635 ;
        RECT 1.510 2.205 2.255 2.375 ;
        RECT 0.085 1.865 1.915 2.035 ;
        RECT 0.085 0.825 0.255 1.865 ;
        RECT 0.990 1.525 1.575 1.695 ;
        RECT 1.405 1.245 1.575 1.525 ;
        RECT 1.745 1.585 1.915 1.865 ;
        RECT 2.085 1.955 2.255 2.205 ;
        RECT 2.085 1.785 3.120 1.955 ;
        RECT 3.290 1.835 3.570 2.635 ;
        RECT 2.950 1.665 3.120 1.785 ;
        RECT 1.745 1.415 2.395 1.585 ;
        RECT 2.950 1.495 3.610 1.665 ;
        RECT 1.405 1.075 1.830 1.245 ;
        RECT 1.405 0.825 1.575 1.075 ;
        RECT 2.225 0.995 2.395 1.415 ;
        RECT 3.440 1.325 3.610 1.495 ;
        RECT 3.440 0.995 3.715 1.325 ;
        RECT 3.440 0.825 3.610 0.995 ;
        RECT 0.085 0.450 0.400 0.825 ;
        RECT 0.655 0.085 0.825 0.825 ;
        RECT 1.075 0.655 1.575 0.825 ;
        RECT 2.015 0.655 3.610 0.825 ;
        RECT 1.075 0.450 1.245 0.655 ;
        RECT 1.470 0.085 1.845 0.485 ;
        RECT 2.015 0.305 2.185 0.655 ;
        RECT 2.370 0.085 2.700 0.485 ;
        RECT 2.870 0.305 3.040 0.655 ;
        RECT 3.210 0.085 3.590 0.485 ;
        RECT 0.000 -0.085 4.140 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
  END
END sky130_fd_sc_hd__or4bb_1

#--------EOF---------

MACRO sky130_fd_sc_hd__or4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4bb_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.640 0.995 3.295 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 2.505 2.125 3.145 2.455 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.430 0.995 0.780 1.695 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.950 0.995 1.240 1.325 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.045 0.785 1.420 1.015 ;
        RECT 3.210 0.785 4.590 1.015 ;
        RECT 0.045 0.335 4.590 0.785 ;
        RECT 0.150 -0.085 0.320 0.335 ;
        RECT 1.430 0.105 4.590 0.335 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.790 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 3.805 1.495 4.080 2.465 ;
        RECT 3.910 0.760 4.080 1.495 ;
        RECT 3.805 0.415 4.080 0.760 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 4.600 2.805 ;
        RECT 0.085 2.035 0.345 2.455 ;
        RECT 0.515 2.205 0.845 2.635 ;
        RECT 1.535 2.205 2.280 2.375 ;
        RECT 0.085 1.865 1.940 2.035 ;
        RECT 0.085 0.825 0.260 1.865 ;
        RECT 0.995 1.525 1.600 1.695 ;
        RECT 1.410 1.245 1.600 1.525 ;
        RECT 1.770 1.585 1.940 1.865 ;
        RECT 2.110 1.955 2.280 2.205 ;
        RECT 2.110 1.785 3.145 1.955 ;
        RECT 3.315 1.835 3.595 2.635 ;
        RECT 2.975 1.665 3.145 1.785 ;
        RECT 1.770 1.415 2.420 1.585 ;
        RECT 2.975 1.495 3.635 1.665 ;
        RECT 1.410 1.075 1.855 1.245 ;
        RECT 1.410 0.825 1.600 1.075 ;
        RECT 2.250 0.995 2.420 1.415 ;
        RECT 3.465 1.325 3.635 1.495 ;
        RECT 4.250 1.440 4.420 2.635 ;
        RECT 3.465 0.995 3.740 1.325 ;
        RECT 3.465 0.825 3.635 0.995 ;
        RECT 0.085 0.450 0.405 0.825 ;
        RECT 0.660 0.085 0.830 0.825 ;
        RECT 1.080 0.655 1.600 0.825 ;
        RECT 2.025 0.655 3.635 0.825 ;
        RECT 1.080 0.450 1.250 0.655 ;
        RECT 1.495 0.085 1.850 0.485 ;
        RECT 2.025 0.305 2.195 0.655 ;
        RECT 2.395 0.085 2.725 0.485 ;
        RECT 2.895 0.305 3.065 0.655 ;
        RECT 3.235 0.085 3.615 0.485 ;
        RECT 4.250 0.085 4.420 1.025 ;
        RECT 0.000 -0.085 4.600 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
  END
END sky130_fd_sc_hd__or4bb_2

#--------EOF---------

MACRO sky130_fd_sc_hd__or4bb_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__or4bb_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 3.235 1.445 3.670 1.615 ;
        RECT 3.235 0.995 3.405 1.445 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 2.795 1.785 3.115 2.375 ;
        RECT 2.795 1.450 3.005 1.785 ;
        RECT 2.675 0.995 3.005 1.450 ;
    END
  END B
  PIN C_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 0.995 0.775 1.695 ;
    END
  END C_N
  PIN D_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 0.945 0.995 1.235 1.325 ;
    END
  END D_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.040 0.335 5.515 1.015 ;
        RECT 0.145 -0.085 0.315 0.335 ;
        RECT 1.425 0.105 5.515 0.335 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 3.875 1.625 4.125 2.465 ;
        RECT 4.715 1.625 4.965 2.465 ;
        RECT 3.875 1.455 5.435 1.625 ;
        RECT 5.205 0.905 5.435 1.455 ;
        RECT 3.915 0.725 5.435 0.905 ;
        RECT 3.915 0.255 4.165 0.725 ;
        RECT 4.675 0.255 5.005 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.085 2.035 0.345 2.455 ;
        RECT 0.515 2.205 0.845 2.635 ;
        RECT 1.125 2.295 2.445 2.465 ;
        RECT 1.125 2.035 1.295 2.295 ;
        RECT 0.085 1.865 1.295 2.035 ;
        RECT 1.510 1.955 2.105 2.125 ;
        RECT 0.085 0.825 0.255 1.865 ;
        RECT 0.990 1.525 1.595 1.695 ;
        RECT 1.405 1.325 1.595 1.525 ;
        RECT 1.405 0.995 1.695 1.325 ;
        RECT 1.405 0.825 1.595 0.995 ;
        RECT 0.085 0.450 0.400 0.825 ;
        RECT 0.655 0.085 0.825 0.825 ;
        RECT 1.075 0.655 1.595 0.825 ;
        RECT 1.935 0.825 2.105 1.955 ;
        RECT 2.275 0.995 2.445 2.295 ;
        RECT 3.400 1.795 3.650 2.635 ;
        RECT 4.295 1.795 4.545 2.635 ;
        RECT 5.135 1.795 5.385 2.635 ;
        RECT 3.575 1.075 5.035 1.245 ;
        RECT 3.575 0.825 3.745 1.075 ;
        RECT 1.935 0.655 3.745 0.825 ;
        RECT 1.075 0.450 1.245 0.655 ;
        RECT 1.515 0.085 1.845 0.480 ;
        RECT 2.095 0.305 2.265 0.655 ;
        RECT 2.465 0.085 2.795 0.485 ;
        RECT 2.965 0.305 3.135 0.655 ;
        RECT 3.355 0.085 3.735 0.485 ;
        RECT 4.335 0.085 4.505 0.555 ;
        RECT 5.175 0.085 5.345 0.555 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
  END
END sky130_fd_sc_hd__or4bb_4

#--------EOF---------

MACRO sky130_fd_sc_hd__probe_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__probe_p_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 1.075 1.240 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.520 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.135 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.520 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 1.250 1.950 4.270 2.160 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.250 0.560 4.270 1.945 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.370 0.680 4.150 1.860 ;
      LAYER via4 ;
        RECT 2.970 0.680 4.150 1.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.395 1.025 4.175 1.355 ;
      LAYER via3 ;
        RECT 3.425 1.030 3.745 1.350 ;
        RECT 3.825 1.030 4.145 1.350 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.095 1.615 0.425 2.465 ;
        RECT 0.595 1.835 0.765 2.635 ;
        RECT 0.935 1.615 1.265 2.465 ;
        RECT 1.435 1.835 1.605 2.635 ;
        RECT 1.855 1.615 2.025 2.465 ;
        RECT 2.195 1.835 2.525 2.635 ;
        RECT 2.695 1.615 2.865 2.465 ;
        RECT 3.035 1.835 3.365 2.635 ;
        RECT 3.535 1.615 3.705 2.465 ;
        RECT 3.875 1.835 4.205 2.635 ;
        RECT 4.375 1.615 4.545 2.465 ;
        RECT 0.095 1.445 1.595 1.615 ;
        RECT 1.855 1.445 4.545 1.615 ;
        RECT 4.715 1.485 5.045 2.635 ;
        RECT 1.420 1.245 1.595 1.445 ;
        RECT 4.290 1.315 4.545 1.445 ;
        RECT 1.420 1.075 4.045 1.245 ;
        RECT 1.420 0.905 1.595 1.075 ;
        RECT 4.290 1.055 4.885 1.315 ;
        RECT 4.290 0.905 4.545 1.055 ;
        RECT 0.175 0.735 1.595 0.905 ;
        RECT 1.855 0.735 4.545 0.905 ;
        RECT 0.175 0.255 0.345 0.735 ;
        RECT 0.515 0.085 0.845 0.565 ;
        RECT 1.015 0.260 1.185 0.735 ;
        RECT 1.355 0.085 1.685 0.565 ;
        RECT 1.855 0.255 2.025 0.735 ;
        RECT 2.195 0.085 2.525 0.565 ;
        RECT 2.695 0.255 2.865 0.735 ;
        RECT 3.035 0.085 3.365 0.565 ;
        RECT 3.535 0.255 3.705 0.735 ;
        RECT 3.875 0.085 4.205 0.565 ;
        RECT 4.375 0.255 4.545 0.735 ;
        RECT 4.715 0.085 5.045 0.885 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 4.320 1.105 4.490 1.275 ;
        RECT 4.680 1.105 4.850 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
      LAYER met1 ;
        RECT 3.465 1.305 4.105 1.320 ;
        RECT 3.465 1.075 4.910 1.305 ;
        RECT 3.465 1.060 4.105 1.075 ;
      LAYER via ;
        RECT 3.495 1.060 3.755 1.320 ;
        RECT 3.815 1.060 4.075 1.320 ;
      LAYER met2 ;
        RECT 3.445 1.005 4.125 1.375 ;
      LAYER via2 ;
        RECT 3.445 1.050 3.725 1.330 ;
        RECT 3.845 1.050 4.125 1.330 ;
  END
END sky130_fd_sc_hd__probe_p_8

#--------EOF---------

MACRO sky130_fd_sc_hd__probec_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__probec_p_8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 1.075 1.240 1.275 ;
    END
  END A
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met5 ;
        RECT 4.360 -0.155 6.675 0.560 ;
        RECT 4.560 -0.455 6.675 -0.155 ;
        RECT 4.360 -1.170 6.675 -0.455 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.930 -0.895 6.110 0.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.130 -0.165 5.910 0.165 ;
      LAYER via3 ;
        RECT 5.160 -0.160 5.480 0.160 ;
        RECT 5.560 -0.160 5.880 0.160 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.135 1.015 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.710 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met5 ;
        RECT 4.360 3.175 6.675 3.890 ;
        RECT 4.560 2.875 6.675 3.175 ;
        RECT 4.360 2.160 6.675 2.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.930 2.435 6.110 3.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.130 2.555 5.910 2.885 ;
      LAYER via3 ;
        RECT 5.160 2.560 5.480 2.880 ;
        RECT 5.560 2.560 5.880 2.880 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT -1.260 0.560 1.060 2.160 ;
    END
    PORT
      LAYER met5 ;
        RECT 1.160 -1.105 2.760 3.825 ;
    END
    PORT
      LAYER met4 ;
        RECT 1.460 0.770 2.640 1.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.885 1.025 2.665 1.355 ;
      LAYER via3 ;
        RECT 1.915 1.030 2.235 1.350 ;
        RECT 2.315 1.030 2.635 1.350 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.890 1.050 2.660 1.330 ;
      LAYER via2 ;
        RECT 1.935 1.050 2.215 1.330 ;
        RECT 2.335 1.050 2.615 1.330 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.520 2.805 ;
        RECT 0.095 1.615 0.425 2.465 ;
        RECT 0.595 1.835 0.765 2.635 ;
        RECT 0.935 1.615 1.265 2.465 ;
        RECT 1.435 1.835 1.605 2.635 ;
        RECT 1.855 1.615 2.025 2.465 ;
        RECT 2.195 1.835 2.525 2.635 ;
        RECT 2.695 1.615 2.865 2.465 ;
        RECT 3.035 1.835 3.365 2.635 ;
        RECT 3.535 1.615 3.705 2.465 ;
        RECT 3.875 1.835 4.205 2.635 ;
        RECT 4.375 1.615 4.545 2.465 ;
        RECT 0.095 1.445 1.595 1.615 ;
        RECT 1.855 1.445 4.545 1.615 ;
        RECT 4.715 1.485 5.045 2.635 ;
        RECT 1.420 1.245 1.595 1.445 ;
        RECT 4.290 1.315 4.545 1.445 ;
        RECT 1.420 1.075 4.045 1.245 ;
        RECT 1.420 0.905 1.595 1.075 ;
        RECT 4.290 1.055 4.870 1.315 ;
        RECT 4.290 0.905 4.545 1.055 ;
        RECT 0.175 0.735 1.595 0.905 ;
        RECT 1.855 0.735 4.545 0.905 ;
        RECT 0.175 0.255 0.345 0.735 ;
        RECT 0.515 0.085 0.845 0.565 ;
        RECT 1.015 0.260 1.185 0.735 ;
        RECT 1.355 0.085 1.685 0.565 ;
        RECT 1.855 0.255 2.025 0.735 ;
        RECT 2.195 0.085 2.525 0.565 ;
        RECT 2.695 0.255 2.865 0.735 ;
        RECT 3.035 0.085 3.365 0.565 ;
        RECT 3.535 0.255 3.705 0.735 ;
        RECT 3.875 0.085 4.205 0.565 ;
        RECT 4.375 0.255 4.545 0.735 ;
        RECT 4.715 0.085 5.045 0.885 ;
        RECT 0.000 -0.085 5.520 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 4.305 1.105 4.475 1.275 ;
        RECT 4.665 1.105 4.835 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
      LAYER met1 ;
        RECT 0.000 2.850 5.520 2.960 ;
        RECT 0.000 2.590 5.840 2.850 ;
        RECT 0.000 2.480 5.520 2.590 ;
        RECT 2.020 1.260 2.660 1.320 ;
        RECT 4.245 1.260 4.895 1.305 ;
        RECT 2.020 1.120 4.895 1.260 ;
        RECT 2.020 1.060 2.660 1.120 ;
        RECT 4.245 1.075 4.895 1.120 ;
        RECT 0.000 0.130 5.520 0.240 ;
        RECT 0.000 -0.130 5.840 0.130 ;
        RECT 0.000 -0.240 5.520 -0.130 ;
      LAYER via ;
        RECT 5.230 2.590 5.490 2.850 ;
        RECT 5.550 2.590 5.810 2.850 ;
        RECT 2.050 1.060 2.310 1.320 ;
        RECT 2.370 1.060 2.630 1.320 ;
        RECT 5.230 -0.130 5.490 0.130 ;
        RECT 5.550 -0.130 5.810 0.130 ;
      LAYER met2 ;
        RECT 5.135 2.580 5.905 2.860 ;
        RECT 5.135 -0.140 5.905 0.140 ;
      LAYER via2 ;
        RECT 5.180 2.580 5.460 2.860 ;
        RECT 5.580 2.580 5.860 2.860 ;
        RECT 5.180 -0.140 5.460 0.140 ;
        RECT 5.580 -0.140 5.860 0.140 ;
      LAYER met3 ;
        RECT -0.715 1.030 0.065 1.350 ;
      LAYER via3 ;
        RECT -0.685 1.030 -0.365 1.350 ;
        RECT -0.285 1.030 0.035 1.350 ;
      LAYER met4 ;
        RECT -1.140 0.770 0.040 1.950 ;
      LAYER met5 ;
        RECT 4.360 2.975 4.460 3.075 ;
        RECT 4.360 -0.355 4.460 -0.255 ;
  END
END sky130_fd_sc_hd__probec_p_8

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfbbn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfbbn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.260 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK_N
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 3.825 1.675 4.060 2.375 ;
        RECT 3.775 1.575 4.060 1.675 ;
        RECT 3.775 1.405 4.105 1.575 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 11.535 1.095 11.990 1.325 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.415 1.025 1.695 1.685 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT 1.935 1.150 2.155 1.695 ;
        RECT 1.935 0.815 2.315 1.150 ;
        RECT 1.935 0.345 2.155 0.815 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 6.065 0.920 6.355 0.965 ;
        RECT 9.745 0.920 10.035 0.965 ;
        RECT 6.065 0.780 10.035 0.920 ;
        RECT 6.065 0.735 6.355 0.780 ;
        RECT 9.745 0.735 10.035 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 14.260 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 11.910 1.005 14.255 1.015 ;
        RECT 6.180 0.785 8.450 1.005 ;
        RECT 10.075 0.785 14.255 1.005 ;
        RECT 0.005 0.105 14.255 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 14.450 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 14.260 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 13.915 1.470 14.175 2.465 ;
        RECT 13.965 0.785 14.175 1.470 ;
        RECT 13.915 0.255 14.175 0.785 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 12.500 1.630 12.785 2.465 ;
        RECT 12.605 0.715 12.785 1.630 ;
        RECT 12.500 0.255 12.785 0.715 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 14.260 2.805 ;
        RECT 0.095 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.095 1.795 0.835 1.965 ;
        RECT 0.605 0.805 0.835 1.795 ;
        RECT 0.095 0.635 0.835 0.805 ;
        RECT 0.095 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.235 2.465 ;
        RECT 1.430 1.885 1.785 2.635 ;
        RECT 2.215 1.875 2.575 2.385 ;
        RECT 2.970 1.905 3.140 2.465 ;
        RECT 3.310 2.215 3.640 2.635 ;
        RECT 4.230 2.135 4.445 2.465 ;
        RECT 4.635 2.250 5.465 2.420 ;
        RECT 2.405 1.505 2.575 1.875 ;
        RECT 2.760 1.745 3.140 1.905 ;
        RECT 2.760 1.575 3.605 1.745 ;
        RECT 2.405 1.465 2.605 1.505 ;
        RECT 2.405 1.430 2.630 1.465 ;
        RECT 2.405 1.405 2.670 1.430 ;
        RECT 2.405 1.295 3.075 1.405 ;
        RECT 2.460 1.255 3.075 1.295 ;
        RECT 2.485 1.075 3.075 1.255 ;
        RECT 3.430 1.095 3.605 1.575 ;
        RECT 4.275 1.305 4.445 2.135 ;
        RECT 4.245 1.275 4.445 1.305 ;
        RECT 4.225 1.235 4.445 1.275 ;
        RECT 3.950 1.175 4.445 1.235 ;
        RECT 4.615 1.575 5.125 1.955 ;
        RECT 3.950 1.105 4.410 1.175 ;
        RECT 1.430 0.085 1.705 0.635 ;
        RECT 2.485 0.595 2.655 1.075 ;
        RECT 3.430 0.795 3.770 1.095 ;
        RECT 2.325 0.265 2.655 0.595 ;
        RECT 2.870 0.765 3.770 0.795 ;
        RECT 3.950 1.065 4.400 1.105 ;
        RECT 2.870 0.625 3.645 0.765 ;
        RECT 2.870 0.305 3.040 0.625 ;
        RECT 3.950 0.595 4.120 1.065 ;
        RECT 4.615 1.035 4.790 1.575 ;
        RECT 5.295 1.405 5.465 2.250 ;
        RECT 5.705 2.205 6.085 2.635 ;
        RECT 6.385 2.035 6.555 2.375 ;
        RECT 5.635 1.785 6.985 2.035 ;
        RECT 7.175 1.915 7.505 2.635 ;
        RECT 8.550 2.250 9.380 2.420 ;
        RECT 9.620 2.255 10.000 2.635 ;
        RECT 5.635 1.575 5.885 1.785 ;
        RECT 6.395 1.405 6.645 1.485 ;
        RECT 5.295 1.235 6.645 1.405 ;
        RECT 5.295 1.195 5.670 1.235 ;
        RECT 4.570 0.705 4.790 1.035 ;
        RECT 5.000 0.735 5.330 1.015 ;
        RECT 5.500 0.655 5.670 1.195 ;
        RECT 6.425 1.155 6.645 1.235 ;
        RECT 6.815 1.065 6.985 1.785 ;
        RECT 7.155 1.415 8.160 1.655 ;
        RECT 8.360 1.575 8.595 1.985 ;
        RECT 7.155 1.235 7.485 1.415 ;
        RECT 8.835 1.305 9.040 1.905 ;
        RECT 7.795 1.065 8.125 1.235 ;
        RECT 5.870 0.965 6.215 1.065 ;
        RECT 6.815 1.060 8.125 1.065 ;
        RECT 5.870 0.735 6.295 0.965 ;
        RECT 6.810 0.895 8.125 1.060 ;
        RECT 8.420 1.125 9.040 1.305 ;
        RECT 9.210 1.405 9.380 2.250 ;
        RECT 10.240 2.085 10.410 2.375 ;
        RECT 10.940 2.255 12.330 2.635 ;
        RECT 9.550 1.915 12.330 2.085 ;
        RECT 9.550 1.575 9.800 1.915 ;
        RECT 9.210 1.235 10.560 1.405 ;
        RECT 6.810 0.780 7.010 0.895 ;
        RECT 3.225 0.085 3.555 0.445 ;
        RECT 3.950 0.425 4.330 0.595 ;
        RECT 5.485 0.585 5.670 0.655 ;
        RECT 6.680 0.610 7.010 0.780 ;
        RECT 5.485 0.465 5.655 0.585 ;
        RECT 4.160 0.265 4.330 0.425 ;
        RECT 4.555 0.265 5.655 0.465 ;
        RECT 5.835 0.085 6.005 0.525 ;
        RECT 6.260 0.425 6.590 0.465 ;
        RECT 7.180 0.425 7.350 0.715 ;
        RECT 8.420 0.705 8.705 1.125 ;
        RECT 9.210 0.465 9.380 1.235 ;
        RECT 10.340 1.075 10.560 1.235 ;
        RECT 9.755 0.735 10.130 1.065 ;
        RECT 10.730 0.780 10.905 1.915 ;
        RECT 10.575 0.595 10.905 0.780 ;
        RECT 11.080 1.575 11.855 1.745 ;
        RECT 11.080 0.925 11.355 1.575 ;
        RECT 12.160 1.325 12.330 1.915 ;
        RECT 12.960 1.325 13.275 2.415 ;
        RECT 13.455 1.765 13.740 2.635 ;
        RECT 12.160 0.995 12.425 1.325 ;
        RECT 12.960 0.995 13.795 1.325 ;
        RECT 11.080 0.755 11.775 0.925 ;
        RECT 6.260 0.255 7.350 0.425 ;
        RECT 7.620 0.085 7.975 0.465 ;
        RECT 8.615 0.265 9.380 0.465 ;
        RECT 9.560 0.085 9.820 0.525 ;
        RECT 10.080 0.425 10.410 0.545 ;
        RECT 11.075 0.425 11.250 0.585 ;
        RECT 10.080 0.255 11.250 0.425 ;
        RECT 11.565 0.265 11.775 0.755 ;
        RECT 12.000 0.085 12.330 0.805 ;
        RECT 12.960 0.255 13.275 0.995 ;
        RECT 13.455 0.085 13.745 0.545 ;
        RECT 0.000 -0.085 14.260 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 0.605 0.765 0.775 0.935 ;
        RECT 1.065 1.785 1.235 1.955 ;
        RECT 2.905 1.105 3.075 1.275 ;
        RECT 4.230 1.105 4.400 1.275 ;
        RECT 4.745 1.785 4.915 1.955 ;
        RECT 5.155 0.765 5.325 0.935 ;
        RECT 8.425 1.785 8.595 1.955 ;
        RECT 7.965 1.445 8.135 1.615 ;
        RECT 6.125 0.765 6.295 0.935 ;
        RECT 8.425 1.105 8.595 1.275 ;
        RECT 9.805 0.765 9.975 0.935 ;
        RECT 11.185 1.445 11.355 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
      LAYER met1 ;
        RECT 1.005 1.940 1.295 1.985 ;
        RECT 4.685 1.940 4.975 1.985 ;
        RECT 8.365 1.940 8.655 1.985 ;
        RECT 1.005 1.800 8.655 1.940 ;
        RECT 1.005 1.755 1.295 1.800 ;
        RECT 4.685 1.755 4.975 1.800 ;
        RECT 8.365 1.755 8.655 1.800 ;
        RECT 7.905 1.600 8.195 1.645 ;
        RECT 11.125 1.600 11.415 1.645 ;
        RECT 7.905 1.460 11.415 1.600 ;
        RECT 7.905 1.415 8.195 1.460 ;
        RECT 11.125 1.415 11.415 1.460 ;
        RECT 2.845 1.260 3.135 1.305 ;
        RECT 4.170 1.260 4.460 1.305 ;
        RECT 8.365 1.260 8.655 1.305 ;
        RECT 2.845 1.120 4.460 1.260 ;
        RECT 2.845 1.075 3.135 1.120 ;
        RECT 4.170 1.075 4.460 1.120 ;
        RECT 5.170 1.120 8.655 1.260 ;
        RECT 5.170 0.965 5.385 1.120 ;
        RECT 8.365 1.075 8.655 1.120 ;
        RECT 0.545 0.920 0.835 0.965 ;
        RECT 5.095 0.920 5.385 0.965 ;
        RECT 0.545 0.780 5.385 0.920 ;
        RECT 0.545 0.735 0.835 0.780 ;
        RECT 5.095 0.735 5.385 0.780 ;
  END
END sky130_fd_sc_hd__sdfbbn_1

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfbbn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfbbn_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.180 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK_N
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 3.825 1.325 4.025 2.375 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 11.590 1.095 12.070 1.325 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.415 1.025 1.695 1.685 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT 1.935 1.095 2.155 1.695 ;
        RECT 1.935 0.765 2.335 1.095 ;
        RECT 1.935 0.345 2.145 0.765 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 6.065 0.920 6.355 0.965 ;
        RECT 9.745 0.920 10.035 0.965 ;
        RECT 6.065 0.780 10.035 0.920 ;
        RECT 6.065 0.735 6.355 0.780 ;
        RECT 9.745 0.735 10.035 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 15.180 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 11.990 1.005 15.175 1.015 ;
        RECT 6.205 0.785 8.475 1.005 ;
        RECT 10.080 0.785 15.175 1.005 ;
        RECT 0.005 0.105 15.175 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 15.370 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 15.180 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 14.415 1.445 14.665 2.465 ;
        RECT 14.460 0.825 14.665 1.445 ;
        RECT 14.415 0.255 14.665 0.825 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 12.580 1.630 12.830 2.465 ;
        RECT 12.660 0.715 12.830 1.630 ;
        RECT 12.580 0.255 12.830 0.715 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 15.180 2.805 ;
        RECT 0.170 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.170 1.795 0.835 1.965 ;
        RECT 0.605 0.805 0.835 1.795 ;
        RECT 0.170 0.635 0.835 0.805 ;
        RECT 0.170 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.235 2.465 ;
        RECT 1.430 1.885 1.785 2.635 ;
        RECT 2.215 1.875 2.575 2.385 ;
        RECT 2.895 1.905 3.065 2.465 ;
        RECT 3.295 2.215 3.640 2.635 ;
        RECT 2.405 1.405 2.575 1.875 ;
        RECT 2.745 1.745 3.065 1.905 ;
        RECT 2.745 1.575 3.645 1.745 ;
        RECT 2.405 1.250 3.075 1.405 ;
        RECT 2.435 1.235 3.075 1.250 ;
        RECT 2.560 1.075 3.075 1.235 ;
        RECT 3.475 1.095 3.645 1.575 ;
        RECT 1.430 0.085 1.705 0.635 ;
        RECT 2.560 0.595 2.730 1.075 ;
        RECT 3.475 0.795 3.770 1.095 ;
        RECT 2.315 0.265 2.730 0.595 ;
        RECT 2.955 0.765 3.770 0.795 ;
        RECT 2.955 0.625 3.645 0.765 ;
        RECT 2.955 0.305 3.125 0.625 ;
        RECT 3.370 0.085 3.700 0.445 ;
        RECT 4.230 0.305 4.455 2.465 ;
        RECT 4.635 2.250 5.465 2.420 ;
        RECT 4.625 1.575 5.125 1.955 ;
        RECT 4.625 0.705 4.845 1.575 ;
        RECT 5.295 1.405 5.465 2.250 ;
        RECT 5.705 2.205 6.085 2.635 ;
        RECT 6.385 2.035 6.555 2.375 ;
        RECT 5.635 1.785 6.985 2.035 ;
        RECT 7.175 1.915 7.505 2.635 ;
        RECT 8.550 2.250 9.380 2.420 ;
        RECT 9.620 2.255 10.000 2.635 ;
        RECT 5.635 1.575 5.885 1.785 ;
        RECT 6.395 1.405 6.645 1.485 ;
        RECT 5.295 1.235 6.645 1.405 ;
        RECT 5.295 1.195 5.715 1.235 ;
        RECT 5.025 0.645 5.375 1.015 ;
        RECT 5.545 0.465 5.715 1.195 ;
        RECT 6.425 1.155 6.645 1.235 ;
        RECT 6.815 1.065 6.985 1.785 ;
        RECT 7.155 1.415 8.160 1.655 ;
        RECT 8.360 1.575 8.595 1.985 ;
        RECT 7.155 1.235 7.485 1.415 ;
        RECT 8.835 1.305 9.040 1.905 ;
        RECT 7.795 1.065 8.125 1.235 ;
        RECT 5.885 0.965 6.215 1.065 ;
        RECT 5.885 0.735 6.295 0.965 ;
        RECT 6.815 0.895 8.125 1.065 ;
        RECT 8.420 1.125 9.040 1.305 ;
        RECT 9.210 1.405 9.380 2.250 ;
        RECT 10.240 2.085 10.410 2.375 ;
        RECT 10.940 2.255 12.410 2.635 ;
        RECT 9.550 1.915 12.410 2.085 ;
        RECT 9.550 1.575 9.800 1.915 ;
        RECT 9.210 1.235 10.560 1.405 ;
        RECT 6.815 0.765 7.035 0.895 ;
        RECT 6.705 0.595 7.035 0.765 ;
        RECT 4.700 0.265 5.715 0.465 ;
        RECT 5.885 0.085 6.055 0.525 ;
        RECT 6.225 0.425 6.555 0.505 ;
        RECT 7.205 0.425 7.375 0.715 ;
        RECT 8.420 0.705 8.705 1.125 ;
        RECT 9.210 0.465 9.380 1.235 ;
        RECT 10.340 1.075 10.560 1.235 ;
        RECT 9.755 0.735 10.130 1.065 ;
        RECT 10.730 0.780 10.910 1.915 ;
        RECT 10.580 0.595 10.910 0.780 ;
        RECT 11.080 1.575 11.925 1.745 ;
        RECT 11.080 0.925 11.355 1.575 ;
        RECT 12.240 1.325 12.410 1.915 ;
        RECT 13.000 1.495 13.235 2.635 ;
        RECT 13.455 1.325 13.770 2.415 ;
        RECT 13.950 1.765 14.245 2.635 ;
        RECT 14.835 1.495 15.075 2.635 ;
        RECT 12.240 0.995 12.480 1.325 ;
        RECT 13.455 0.995 14.290 1.325 ;
        RECT 11.080 0.755 11.845 0.925 ;
        RECT 6.225 0.255 7.375 0.425 ;
        RECT 7.645 0.085 7.975 0.465 ;
        RECT 8.615 0.265 9.380 0.465 ;
        RECT 9.560 0.085 9.820 0.525 ;
        RECT 10.080 0.425 10.410 0.545 ;
        RECT 11.080 0.425 11.250 0.585 ;
        RECT 10.080 0.255 11.250 0.425 ;
        RECT 11.620 0.265 11.845 0.755 ;
        RECT 12.080 0.085 12.410 0.805 ;
        RECT 13.000 0.085 13.235 0.885 ;
        RECT 13.455 0.255 13.770 0.995 ;
        RECT 13.950 0.085 14.245 0.545 ;
        RECT 14.835 0.085 15.075 0.885 ;
        RECT 0.000 -0.085 15.180 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 0.605 0.765 0.775 0.935 ;
        RECT 1.065 1.785 1.235 1.955 ;
        RECT 2.905 1.105 3.075 1.275 ;
        RECT 4.285 1.105 4.455 1.275 ;
        RECT 4.745 1.785 4.915 1.955 ;
        RECT 5.205 0.765 5.375 0.935 ;
        RECT 8.425 1.785 8.595 1.955 ;
        RECT 7.965 1.445 8.135 1.615 ;
        RECT 6.125 0.765 6.295 0.935 ;
        RECT 8.425 1.105 8.595 1.275 ;
        RECT 9.805 0.765 9.975 0.935 ;
        RECT 11.185 1.445 11.355 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
      LAYER met1 ;
        RECT 1.005 1.940 1.295 1.985 ;
        RECT 4.685 1.940 4.975 1.985 ;
        RECT 8.365 1.940 8.655 1.985 ;
        RECT 1.005 1.800 8.655 1.940 ;
        RECT 1.005 1.755 1.295 1.800 ;
        RECT 4.685 1.755 4.975 1.800 ;
        RECT 8.365 1.755 8.655 1.800 ;
        RECT 7.905 1.600 8.195 1.645 ;
        RECT 11.125 1.600 11.415 1.645 ;
        RECT 7.905 1.460 11.415 1.600 ;
        RECT 7.905 1.415 8.195 1.460 ;
        RECT 11.125 1.415 11.415 1.460 ;
        RECT 2.845 1.260 3.135 1.305 ;
        RECT 4.225 1.260 4.515 1.305 ;
        RECT 8.365 1.260 8.655 1.305 ;
        RECT 2.845 1.120 4.515 1.260 ;
        RECT 2.845 1.075 3.135 1.120 ;
        RECT 4.225 1.075 4.515 1.120 ;
        RECT 5.220 1.120 8.655 1.260 ;
        RECT 5.220 0.965 5.435 1.120 ;
        RECT 8.365 1.075 8.655 1.120 ;
        RECT 0.545 0.920 0.835 0.965 ;
        RECT 5.145 0.920 5.435 0.965 ;
        RECT 0.545 0.780 5.435 0.920 ;
        RECT 0.545 0.735 0.835 0.780 ;
        RECT 5.145 0.735 5.435 0.780 ;
  END
END sky130_fd_sc_hd__sdfbbn_2

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfbbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfbbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.260 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.975 0.435 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER li1 ;
        RECT 3.825 1.325 4.025 2.375 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 11.535 1.095 11.990 1.325 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.440 1.025 1.720 1.685 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER li1 ;
        RECT 1.960 1.015 2.180 1.695 ;
        RECT 1.960 0.845 2.415 1.015 ;
        RECT 1.960 0.345 2.180 0.845 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 6.065 0.920 6.355 0.965 ;
        RECT 9.745 0.920 10.035 0.965 ;
        RECT 6.065 0.780 10.035 0.920 ;
        RECT 6.065 0.735 6.355 0.780 ;
        RECT 9.745 0.735 10.035 0.780 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 14.260 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 11.910 1.005 14.255 1.015 ;
        RECT 6.200 0.785 8.470 1.005 ;
        RECT 10.075 0.785 14.255 1.005 ;
        RECT 0.005 0.105 14.255 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 14.450 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 14.260 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 13.915 1.605 14.175 2.465 ;
        RECT 13.965 0.825 14.175 1.605 ;
        RECT 13.915 0.255 14.175 0.825 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 12.500 1.630 12.785 2.465 ;
        RECT 12.605 0.715 12.785 1.630 ;
        RECT 12.500 0.255 12.785 0.715 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 14.260 2.805 ;
        RECT 0.170 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.170 1.795 0.835 1.965 ;
        RECT 0.605 0.805 0.835 1.795 ;
        RECT 0.170 0.635 0.835 0.805 ;
        RECT 0.170 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.240 2.465 ;
        RECT 1.455 1.885 1.785 2.635 ;
        RECT 2.235 1.875 2.565 2.385 ;
        RECT 2.895 1.905 3.065 2.465 ;
        RECT 3.310 2.215 3.640 2.635 ;
        RECT 2.350 1.365 2.565 1.875 ;
        RECT 2.745 1.745 3.065 1.905 ;
        RECT 2.745 1.575 3.645 1.745 ;
        RECT 2.350 1.185 3.075 1.365 ;
        RECT 2.585 1.075 3.075 1.185 ;
        RECT 3.475 1.095 3.645 1.575 ;
        RECT 1.455 0.085 1.705 0.635 ;
        RECT 2.585 0.595 2.755 1.075 ;
        RECT 3.475 0.795 3.770 1.095 ;
        RECT 2.350 0.265 2.755 0.595 ;
        RECT 2.925 0.765 3.770 0.795 ;
        RECT 2.925 0.625 3.645 0.765 ;
        RECT 2.925 0.305 3.125 0.625 ;
        RECT 3.370 0.085 3.700 0.445 ;
        RECT 4.230 0.305 4.455 2.465 ;
        RECT 4.635 2.250 5.465 2.420 ;
        RECT 4.625 1.575 5.125 1.955 ;
        RECT 4.625 0.705 4.845 1.575 ;
        RECT 5.295 1.405 5.465 2.250 ;
        RECT 5.705 2.205 6.085 2.635 ;
        RECT 6.385 2.035 6.555 2.375 ;
        RECT 5.635 1.785 6.985 2.035 ;
        RECT 7.175 1.915 7.505 2.635 ;
        RECT 8.550 2.250 9.380 2.420 ;
        RECT 9.620 2.255 10.000 2.635 ;
        RECT 5.635 1.575 5.885 1.785 ;
        RECT 6.395 1.405 6.645 1.485 ;
        RECT 5.295 1.235 6.645 1.405 ;
        RECT 5.295 1.195 5.715 1.235 ;
        RECT 5.025 0.645 5.375 1.015 ;
        RECT 5.545 0.465 5.715 1.195 ;
        RECT 6.425 1.155 6.645 1.235 ;
        RECT 6.815 1.065 6.985 1.785 ;
        RECT 7.155 1.415 8.160 1.655 ;
        RECT 8.360 1.575 8.595 1.985 ;
        RECT 7.155 1.235 7.485 1.415 ;
        RECT 8.835 1.305 9.040 1.905 ;
        RECT 7.795 1.065 8.125 1.235 ;
        RECT 5.885 0.965 6.215 1.065 ;
        RECT 5.885 0.735 6.295 0.965 ;
        RECT 6.815 0.895 8.125 1.065 ;
        RECT 8.420 1.125 9.040 1.305 ;
        RECT 9.210 1.405 9.380 2.250 ;
        RECT 10.240 2.085 10.410 2.375 ;
        RECT 10.940 2.255 12.330 2.635 ;
        RECT 9.550 1.915 12.330 2.085 ;
        RECT 9.550 1.575 9.800 1.915 ;
        RECT 9.210 1.235 10.560 1.405 ;
        RECT 6.815 0.765 7.030 0.895 ;
        RECT 6.700 0.595 7.030 0.765 ;
        RECT 4.700 0.265 5.715 0.465 ;
        RECT 5.885 0.085 6.055 0.525 ;
        RECT 6.225 0.425 6.555 0.465 ;
        RECT 7.200 0.425 7.395 0.715 ;
        RECT 8.420 0.705 8.705 1.125 ;
        RECT 9.210 0.465 9.380 1.235 ;
        RECT 10.340 1.075 10.560 1.235 ;
        RECT 9.755 0.735 10.130 1.065 ;
        RECT 10.730 0.815 10.905 1.915 ;
        RECT 10.575 0.645 10.905 0.815 ;
        RECT 11.080 1.575 11.855 1.745 ;
        RECT 11.080 0.925 11.355 1.575 ;
        RECT 12.160 1.325 12.330 1.915 ;
        RECT 12.960 1.325 13.275 2.415 ;
        RECT 13.450 1.765 13.745 2.635 ;
        RECT 12.160 0.995 12.425 1.325 ;
        RECT 12.960 0.995 13.795 1.325 ;
        RECT 11.080 0.755 11.765 0.925 ;
        RECT 6.225 0.255 7.395 0.425 ;
        RECT 7.640 0.085 7.975 0.465 ;
        RECT 8.615 0.265 9.380 0.465 ;
        RECT 9.560 0.085 9.820 0.525 ;
        RECT 10.080 0.425 10.430 0.465 ;
        RECT 11.075 0.425 11.250 0.585 ;
        RECT 10.080 0.255 11.250 0.425 ;
        RECT 11.565 0.265 11.765 0.755 ;
        RECT 12.000 0.085 12.330 0.805 ;
        RECT 12.960 0.255 13.275 0.995 ;
        RECT 13.455 0.085 13.745 0.545 ;
        RECT 0.000 -0.085 14.260 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 0.605 1.785 0.775 1.955 ;
        RECT 1.065 0.765 1.235 0.935 ;
        RECT 2.905 1.105 3.075 1.275 ;
        RECT 4.285 1.105 4.455 1.275 ;
        RECT 4.745 1.785 4.915 1.955 ;
        RECT 5.205 0.765 5.375 0.935 ;
        RECT 8.425 1.785 8.595 1.955 ;
        RECT 7.965 1.445 8.135 1.615 ;
        RECT 6.125 0.765 6.295 0.935 ;
        RECT 8.425 1.105 8.595 1.275 ;
        RECT 9.805 0.765 9.975 0.935 ;
        RECT 11.185 1.445 11.355 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
      LAYER met1 ;
        RECT 0.545 1.940 0.835 1.985 ;
        RECT 4.685 1.940 4.975 1.985 ;
        RECT 8.365 1.940 8.655 1.985 ;
        RECT 0.545 1.800 8.655 1.940 ;
        RECT 0.545 1.755 0.835 1.800 ;
        RECT 4.685 1.755 4.975 1.800 ;
        RECT 8.365 1.755 8.655 1.800 ;
        RECT 7.905 1.600 8.195 1.645 ;
        RECT 11.125 1.600 11.415 1.645 ;
        RECT 7.905 1.460 11.415 1.600 ;
        RECT 7.905 1.415 8.195 1.460 ;
        RECT 11.125 1.415 11.415 1.460 ;
        RECT 2.845 1.260 3.135 1.305 ;
        RECT 4.225 1.260 4.515 1.305 ;
        RECT 8.365 1.260 8.655 1.305 ;
        RECT 2.845 1.120 4.515 1.260 ;
        RECT 2.845 1.075 3.135 1.120 ;
        RECT 4.225 1.075 4.515 1.120 ;
        RECT 5.220 1.120 8.655 1.260 ;
        RECT 5.220 0.965 5.435 1.120 ;
        RECT 8.365 1.075 8.655 1.120 ;
        RECT 1.005 0.920 1.295 0.965 ;
        RECT 5.145 0.920 5.435 0.965 ;
        RECT 1.005 0.780 5.435 0.920 ;
        RECT 1.005 0.735 1.295 0.780 ;
        RECT 5.145 0.735 5.435 0.780 ;
  END
END sky130_fd_sc_hd__sdfbbp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.975 0.490 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.144000 ;
    PORT
      LAYER li1 ;
        RECT 2.865 1.785 3.120 2.465 ;
        RECT 2.735 1.355 3.120 1.785 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 9.630 0.965 9.920 1.305 ;
        RECT 6.445 0.920 7.095 0.965 ;
        RECT 9.630 0.920 10.175 0.965 ;
        RECT 6.445 0.780 10.175 0.920 ;
        RECT 6.445 0.735 7.095 0.780 ;
        RECT 9.885 0.735 10.175 0.780 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.156600 ;
    PORT
      LAYER li1 ;
        RECT 4.020 0.710 4.395 1.700 ;
        RECT 4.020 0.285 4.275 0.710 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.730 2.465 ;
        RECT 1.485 1.070 1.730 1.985 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.880 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.880 1.355 1.015 ;
        RECT 2.305 0.880 3.640 1.145 ;
        RECT 0.005 0.725 4.885 0.880 ;
        RECT 6.955 0.785 7.865 1.005 ;
        RECT 10.550 0.885 11.480 1.015 ;
        RECT 10.550 0.785 12.860 0.885 ;
        RECT 5.935 0.725 12.860 0.785 ;
        RECT 0.005 0.465 12.860 0.725 ;
        RECT 0.005 0.200 2.295 0.465 ;
        RECT 3.150 0.200 12.860 0.465 ;
        RECT 0.005 0.105 1.355 0.200 ;
        RECT 4.895 0.105 12.860 0.200 ;
        RECT 0.215 -0.010 0.235 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.425 13.070 2.910 ;
        RECT -0.190 1.305 1.970 1.425 ;
        RECT 4.405 1.305 13.070 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 12.880 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 11.140 1.460 11.400 2.325 ;
        RECT 11.150 1.445 11.400 1.460 ;
        RECT 11.190 0.795 11.400 1.445 ;
        RECT 11.140 0.265 11.400 0.795 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER li1 ;
        RECT 12.510 1.560 12.780 2.465 ;
        RECT 12.600 0.760 12.780 1.560 ;
        RECT 12.520 0.255 12.780 0.760 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 12.880 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.530 2.135 0.860 2.635 ;
        RECT 0.090 1.795 0.865 1.965 ;
        RECT 0.660 1.325 0.865 1.795 ;
        RECT 1.035 1.900 1.205 2.465 ;
        RECT 1.900 2.055 2.150 2.400 ;
        RECT 1.035 1.730 1.315 1.900 ;
        RECT 0.660 0.995 0.975 1.325 ;
        RECT 0.660 0.805 0.835 0.995 ;
        RECT 0.095 0.635 0.835 0.805 ;
        RECT 1.145 0.675 1.315 1.730 ;
        RECT 1.980 1.455 2.150 2.055 ;
        RECT 2.320 2.040 2.490 2.635 ;
        RECT 3.460 2.105 3.630 2.465 ;
        RECT 4.300 2.275 4.630 2.635 ;
        RECT 4.905 2.185 5.275 2.435 ;
        RECT 4.905 2.105 5.075 2.185 ;
        RECT 5.470 2.135 5.835 2.465 ;
        RECT 3.290 1.935 5.075 2.105 ;
        RECT 1.980 1.260 2.470 1.455 ;
        RECT 2.055 1.185 2.470 1.260 ;
        RECT 3.290 1.185 3.460 1.935 ;
        RECT 2.055 0.995 3.085 1.185 ;
        RECT 2.055 0.900 2.225 0.995 ;
        RECT 0.095 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.315 0.675 ;
        RECT 1.535 0.730 2.225 0.900 ;
        RECT 1.535 0.395 1.705 0.730 ;
        RECT 1.875 0.085 2.205 0.560 ;
        RECT 2.395 0.085 2.725 0.825 ;
        RECT 2.915 0.425 3.085 0.995 ;
        RECT 3.255 1.015 3.460 1.185 ;
        RECT 3.255 0.675 3.425 1.015 ;
        RECT 3.680 0.425 3.850 1.685 ;
        RECT 4.565 0.895 4.735 1.935 ;
        RECT 5.245 1.575 5.495 1.955 ;
        RECT 4.905 1.065 5.075 1.395 ;
        RECT 5.325 1.035 5.495 1.575 ;
        RECT 5.665 1.385 5.835 2.135 ;
        RECT 6.005 2.105 6.175 2.375 ;
        RECT 6.410 2.355 6.740 2.635 ;
        RECT 6.995 2.105 7.165 2.375 ;
        RECT 7.375 2.175 7.745 2.635 ;
        RECT 6.005 1.935 7.165 2.105 ;
        RECT 7.970 2.005 8.140 2.465 ;
        RECT 8.320 2.125 9.190 2.465 ;
        RECT 9.360 2.195 9.610 2.635 ;
        RECT 9.015 2.115 9.190 2.125 ;
        RECT 9.015 2.035 9.210 2.115 ;
        RECT 7.455 1.835 8.140 2.005 ;
        RECT 8.310 1.935 8.840 1.955 ;
        RECT 7.455 1.765 7.715 1.835 ;
        RECT 6.285 1.595 7.715 1.765 ;
        RECT 8.310 1.665 8.870 1.935 ;
        RECT 5.665 1.215 7.375 1.385 ;
        RECT 4.565 0.715 5.145 0.895 ;
        RECT 2.915 0.255 3.850 0.425 ;
        RECT 4.445 0.085 4.775 0.540 ;
        RECT 4.975 0.505 5.145 0.715 ;
        RECT 5.325 0.705 5.975 1.035 ;
        RECT 4.975 0.335 5.315 0.505 ;
        RECT 6.165 0.475 6.335 1.215 ;
        RECT 6.505 0.765 7.035 1.045 ;
        RECT 7.205 1.005 7.375 1.215 ;
        RECT 7.545 0.835 7.715 1.595 ;
        RECT 5.485 0.305 6.335 0.475 ;
        RECT 6.915 0.085 7.245 0.545 ;
        RECT 7.455 0.445 7.715 0.835 ;
        RECT 7.885 1.655 8.870 1.665 ;
        RECT 9.040 1.745 9.210 2.035 ;
        RECT 9.780 2.085 9.950 2.375 ;
        RECT 10.120 2.255 10.450 2.635 ;
        RECT 9.780 1.915 10.545 2.085 ;
        RECT 7.885 1.495 8.520 1.655 ;
        RECT 9.040 1.575 10.205 1.745 ;
        RECT 7.885 0.705 8.095 1.495 ;
        RECT 9.040 1.485 9.210 1.575 ;
        RECT 8.405 0.920 8.575 1.325 ;
        RECT 8.745 1.315 9.210 1.485 ;
        RECT 10.375 1.325 10.545 1.915 ;
        RECT 10.720 1.495 10.970 2.635 ;
        RECT 11.650 1.705 11.830 2.465 ;
        RECT 12.010 1.875 12.340 2.635 ;
        RECT 11.650 1.535 12.325 1.705 ;
        RECT 12.155 1.390 12.325 1.535 ;
        RECT 8.745 0.535 8.915 1.315 ;
        RECT 10.375 1.295 11.020 1.325 ;
        RECT 9.125 0.865 9.295 1.145 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.125 0.695 9.655 0.865 ;
        RECT 7.455 0.275 7.785 0.445 ;
        RECT 8.005 0.255 8.915 0.535 ;
        RECT 9.085 0.085 9.255 0.525 ;
        RECT 9.485 0.465 9.655 0.695 ;
        RECT 9.825 0.635 10.115 1.065 ;
        RECT 10.345 0.995 11.020 1.295 ;
        RECT 12.155 1.060 12.430 1.390 ;
        RECT 10.345 0.465 10.515 0.995 ;
        RECT 12.155 0.805 12.325 1.060 ;
        RECT 11.660 0.635 12.325 0.805 ;
        RECT 9.485 0.295 10.515 0.465 ;
        RECT 10.720 0.085 10.890 0.545 ;
        RECT 11.660 0.255 11.830 0.635 ;
        RECT 12.010 0.085 12.340 0.465 ;
        RECT 0.000 -0.085 12.880 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 1.035 1.785 1.205 1.955 ;
        RECT 0.805 1.105 0.975 1.275 ;
        RECT 5.325 1.785 5.495 1.955 ;
        RECT 4.905 1.105 5.075 1.275 ;
        RECT 8.445 1.785 8.615 1.955 ;
        RECT 6.865 0.765 7.035 0.935 ;
        RECT 8.405 1.105 8.575 1.275 ;
        RECT 9.690 1.105 9.860 1.275 ;
        RECT 9.945 0.765 10.115 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
      LAYER met1 ;
        RECT 0.970 1.940 1.270 1.985 ;
        RECT 5.265 1.940 5.555 1.985 ;
        RECT 8.385 1.940 8.675 1.985 ;
        RECT 0.970 1.800 8.675 1.940 ;
        RECT 0.970 1.755 1.270 1.800 ;
        RECT 5.265 1.755 5.555 1.800 ;
        RECT 8.385 1.755 8.675 1.800 ;
        RECT 0.745 1.260 1.035 1.305 ;
        RECT 4.845 1.260 5.135 1.305 ;
        RECT 8.345 1.260 8.635 1.305 ;
        RECT 0.745 1.120 8.635 1.260 ;
        RECT 0.745 1.075 1.035 1.120 ;
        RECT 4.845 1.075 5.135 1.120 ;
        RECT 8.345 1.075 8.635 1.120 ;
  END
END sky130_fd_sc_hd__sdfrbp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.340 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.975 0.490 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.144000 ;
    PORT
      LAYER li1 ;
        RECT 2.865 1.785 3.120 2.465 ;
        RECT 2.735 1.355 3.120 1.785 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 9.630 0.965 9.920 1.305 ;
        RECT 6.445 0.920 7.095 0.965 ;
        RECT 9.630 0.920 10.175 0.965 ;
        RECT 6.445 0.780 10.175 0.920 ;
        RECT 6.445 0.735 7.095 0.780 ;
        RECT 9.885 0.735 10.175 0.780 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.156600 ;
    PORT
      LAYER li1 ;
        RECT 4.020 0.710 4.395 1.700 ;
        RECT 4.020 0.285 4.275 0.710 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.730 2.465 ;
        RECT 1.485 1.070 1.730 1.985 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 13.340 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.880 1.355 1.015 ;
        RECT 2.305 0.880 3.640 1.145 ;
        RECT 0.005 0.725 4.885 0.880 ;
        RECT 6.955 0.785 7.865 1.005 ;
        RECT 11.030 0.785 13.335 1.015 ;
        RECT 5.935 0.725 13.335 0.785 ;
        RECT 0.005 0.465 13.335 0.725 ;
        RECT 0.005 0.200 2.295 0.465 ;
        RECT 3.150 0.200 13.335 0.465 ;
        RECT 0.005 0.105 1.355 0.200 ;
        RECT 4.895 0.105 13.335 0.200 ;
        RECT 0.215 -0.010 0.235 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.425 13.530 2.910 ;
        RECT -0.190 1.305 1.970 1.425 ;
        RECT 4.405 1.305 13.530 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 13.340 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.511500 ;
    PORT
      LAYER li1 ;
        RECT 11.575 0.265 11.925 1.695 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 12.525 2.080 12.825 2.465 ;
        RECT 12.435 1.535 12.825 2.080 ;
        RECT 12.655 0.825 12.825 1.535 ;
        RECT 12.445 0.310 12.825 0.825 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 13.340 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.530 2.135 0.860 2.635 ;
        RECT 0.090 1.795 0.865 1.965 ;
        RECT 0.660 1.325 0.865 1.795 ;
        RECT 1.035 1.900 1.205 2.465 ;
        RECT 1.900 2.055 2.150 2.400 ;
        RECT 1.035 1.730 1.315 1.900 ;
        RECT 0.660 0.995 0.975 1.325 ;
        RECT 0.660 0.805 0.835 0.995 ;
        RECT 0.095 0.635 0.835 0.805 ;
        RECT 1.145 0.675 1.315 1.730 ;
        RECT 1.980 1.455 2.150 2.055 ;
        RECT 2.320 2.040 2.490 2.635 ;
        RECT 3.460 2.105 3.630 2.465 ;
        RECT 4.300 2.275 4.630 2.635 ;
        RECT 4.905 2.185 5.275 2.435 ;
        RECT 4.905 2.105 5.075 2.185 ;
        RECT 5.470 2.135 5.835 2.465 ;
        RECT 3.290 1.935 5.075 2.105 ;
        RECT 1.980 1.260 2.470 1.455 ;
        RECT 2.055 1.185 2.470 1.260 ;
        RECT 3.290 1.185 3.460 1.935 ;
        RECT 2.055 0.995 3.085 1.185 ;
        RECT 2.055 0.900 2.225 0.995 ;
        RECT 0.095 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.315 0.675 ;
        RECT 1.535 0.730 2.225 0.900 ;
        RECT 1.535 0.395 1.705 0.730 ;
        RECT 1.875 0.085 2.205 0.560 ;
        RECT 2.395 0.085 2.725 0.825 ;
        RECT 2.915 0.425 3.085 0.995 ;
        RECT 3.255 1.015 3.460 1.185 ;
        RECT 3.255 0.675 3.425 1.015 ;
        RECT 3.680 0.425 3.850 1.685 ;
        RECT 4.565 0.895 4.735 1.935 ;
        RECT 5.245 1.575 5.495 1.955 ;
        RECT 4.905 1.065 5.075 1.395 ;
        RECT 5.325 1.035 5.495 1.575 ;
        RECT 5.665 1.385 5.835 2.135 ;
        RECT 6.005 2.105 6.175 2.375 ;
        RECT 6.410 2.355 6.740 2.635 ;
        RECT 6.995 2.105 7.165 2.375 ;
        RECT 7.375 2.175 7.745 2.635 ;
        RECT 6.005 1.935 7.165 2.105 ;
        RECT 7.970 2.005 8.140 2.465 ;
        RECT 8.320 2.125 9.190 2.465 ;
        RECT 9.360 2.195 9.610 2.635 ;
        RECT 9.015 2.115 9.190 2.125 ;
        RECT 9.015 2.035 9.210 2.115 ;
        RECT 7.455 1.835 8.140 2.005 ;
        RECT 8.310 1.935 8.840 1.955 ;
        RECT 7.455 1.765 7.715 1.835 ;
        RECT 6.285 1.595 7.715 1.765 ;
        RECT 8.310 1.665 8.870 1.935 ;
        RECT 5.665 1.215 7.375 1.385 ;
        RECT 4.565 0.715 5.145 0.895 ;
        RECT 2.915 0.255 3.850 0.425 ;
        RECT 4.445 0.085 4.775 0.540 ;
        RECT 4.975 0.505 5.145 0.715 ;
        RECT 5.325 0.705 5.975 1.035 ;
        RECT 4.975 0.335 5.315 0.505 ;
        RECT 6.165 0.475 6.335 1.215 ;
        RECT 6.505 0.765 7.035 1.045 ;
        RECT 7.205 1.005 7.375 1.215 ;
        RECT 7.545 0.835 7.715 1.595 ;
        RECT 5.485 0.305 6.335 0.475 ;
        RECT 6.915 0.085 7.245 0.545 ;
        RECT 7.455 0.445 7.715 0.835 ;
        RECT 7.885 1.655 8.870 1.665 ;
        RECT 9.040 1.745 9.210 2.035 ;
        RECT 9.780 2.085 9.950 2.375 ;
        RECT 10.120 2.255 10.450 2.635 ;
        RECT 9.780 1.915 10.545 2.085 ;
        RECT 7.885 1.495 8.520 1.655 ;
        RECT 9.040 1.575 10.205 1.745 ;
        RECT 7.885 0.705 8.095 1.495 ;
        RECT 9.040 1.485 9.210 1.575 ;
        RECT 8.405 0.920 8.575 1.325 ;
        RECT 8.745 1.315 9.210 1.485 ;
        RECT 10.375 1.325 10.545 1.915 ;
        RECT 10.715 2.035 10.890 2.465 ;
        RECT 11.090 2.205 11.420 2.635 ;
        RECT 12.025 2.255 12.355 2.635 ;
        RECT 11.550 2.035 12.265 2.085 ;
        RECT 10.715 1.865 12.265 2.035 ;
        RECT 10.715 1.795 11.405 1.865 ;
        RECT 8.745 0.535 8.915 1.315 ;
        RECT 10.375 1.295 11.060 1.325 ;
        RECT 9.125 0.865 9.295 1.145 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.125 0.695 9.655 0.865 ;
        RECT 7.455 0.275 7.785 0.445 ;
        RECT 8.005 0.255 8.915 0.535 ;
        RECT 9.085 0.085 9.255 0.525 ;
        RECT 9.485 0.465 9.655 0.695 ;
        RECT 9.825 0.635 10.115 1.065 ;
        RECT 10.345 1.055 11.060 1.295 ;
        RECT 10.345 0.465 10.515 1.055 ;
        RECT 11.230 0.885 11.405 1.795 ;
        RECT 12.095 1.325 12.265 1.865 ;
        RECT 12.995 1.495 13.245 2.635 ;
        RECT 12.095 0.995 12.485 1.325 ;
        RECT 9.485 0.295 10.515 0.465 ;
        RECT 10.715 0.715 11.405 0.885 ;
        RECT 10.715 0.345 10.885 0.715 ;
        RECT 11.090 0.085 11.365 0.545 ;
        RECT 12.105 0.085 12.275 0.825 ;
        RECT 12.995 0.085 13.165 0.930 ;
        RECT 0.000 -0.085 13.340 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 1.035 1.785 1.205 1.955 ;
        RECT 0.805 1.105 0.975 1.275 ;
        RECT 5.325 1.785 5.495 1.955 ;
        RECT 4.905 1.105 5.075 1.275 ;
        RECT 8.445 1.785 8.615 1.955 ;
        RECT 6.865 0.765 7.035 0.935 ;
        RECT 8.405 1.105 8.575 1.275 ;
        RECT 9.690 1.105 9.860 1.275 ;
        RECT 9.945 0.765 10.115 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
      LAYER met1 ;
        RECT 0.970 1.940 1.270 1.985 ;
        RECT 5.265 1.940 5.555 1.985 ;
        RECT 8.385 1.940 8.675 1.985 ;
        RECT 0.970 1.800 8.675 1.940 ;
        RECT 0.970 1.755 1.270 1.800 ;
        RECT 5.265 1.755 5.555 1.800 ;
        RECT 8.385 1.755 8.675 1.800 ;
        RECT 0.745 1.260 1.035 1.305 ;
        RECT 4.845 1.260 5.135 1.305 ;
        RECT 8.345 1.260 8.635 1.305 ;
        RECT 0.745 1.120 8.635 1.260 ;
        RECT 0.745 1.075 1.035 1.120 ;
        RECT 4.845 1.075 5.135 1.120 ;
        RECT 8.345 1.075 8.635 1.120 ;
  END
END sky130_fd_sc_hd__sdfrbp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfrtn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtn_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.500 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK_N
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.975 0.490 1.625 ;
    END
  END CLK_N
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.144000 ;
    PORT
      LAYER li1 ;
        RECT 2.865 1.785 3.120 2.465 ;
        RECT 2.735 1.355 3.120 1.785 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 9.630 0.965 9.920 1.305 ;
        RECT 6.445 0.920 7.095 0.965 ;
        RECT 9.630 0.920 10.175 0.965 ;
        RECT 6.445 0.780 10.175 0.920 ;
        RECT 6.445 0.735 7.095 0.780 ;
        RECT 9.885 0.735 10.175 0.780 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.156600 ;
    PORT
      LAYER li1 ;
        RECT 4.020 0.710 4.395 1.700 ;
        RECT 4.020 0.285 4.275 0.710 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.730 2.465 ;
        RECT 1.485 1.070 1.730 1.985 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.500 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.880 1.355 1.015 ;
        RECT 2.305 0.880 3.640 1.145 ;
        RECT 0.005 0.725 4.885 0.880 ;
        RECT 6.955 0.785 7.865 1.005 ;
        RECT 10.550 0.785 11.480 1.015 ;
        RECT 5.935 0.725 11.480 0.785 ;
        RECT 0.005 0.465 11.480 0.725 ;
        RECT 0.005 0.200 2.295 0.465 ;
        RECT 3.150 0.200 11.480 0.465 ;
        RECT 0.005 0.105 1.355 0.200 ;
        RECT 4.895 0.105 11.480 0.200 ;
        RECT 0.215 -0.010 0.235 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.425 11.690 2.910 ;
        RECT -0.190 1.305 1.970 1.425 ;
        RECT 4.405 1.305 11.690 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.500 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 11.140 1.460 11.400 2.325 ;
        RECT 11.150 1.445 11.400 1.460 ;
        RECT 11.190 0.795 11.400 1.445 ;
        RECT 11.140 0.265 11.400 0.795 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.500 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.530 2.135 0.860 2.635 ;
        RECT 0.090 1.795 0.865 1.965 ;
        RECT 0.660 1.325 0.865 1.795 ;
        RECT 1.035 1.900 1.205 2.465 ;
        RECT 1.900 2.055 2.150 2.400 ;
        RECT 1.035 1.730 1.315 1.900 ;
        RECT 0.660 0.995 0.975 1.325 ;
        RECT 0.660 0.805 0.835 0.995 ;
        RECT 0.095 0.635 0.835 0.805 ;
        RECT 1.145 0.675 1.315 1.730 ;
        RECT 1.980 1.455 2.150 2.055 ;
        RECT 2.320 2.040 2.490 2.635 ;
        RECT 3.460 2.105 3.630 2.465 ;
        RECT 4.300 2.275 4.630 2.635 ;
        RECT 4.905 2.185 5.275 2.435 ;
        RECT 4.905 2.105 5.075 2.185 ;
        RECT 5.470 2.135 5.835 2.465 ;
        RECT 3.290 1.935 5.075 2.105 ;
        RECT 1.980 1.260 2.470 1.455 ;
        RECT 2.055 1.185 2.470 1.260 ;
        RECT 3.290 1.185 3.460 1.935 ;
        RECT 2.055 0.995 3.085 1.185 ;
        RECT 2.055 0.900 2.225 0.995 ;
        RECT 0.095 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.315 0.675 ;
        RECT 1.535 0.730 2.225 0.900 ;
        RECT 1.535 0.395 1.705 0.730 ;
        RECT 1.875 0.085 2.205 0.560 ;
        RECT 2.395 0.085 2.725 0.825 ;
        RECT 2.915 0.425 3.085 0.995 ;
        RECT 3.255 1.015 3.460 1.185 ;
        RECT 3.255 0.675 3.425 1.015 ;
        RECT 3.680 0.425 3.850 1.685 ;
        RECT 4.565 0.895 4.735 1.935 ;
        RECT 5.245 1.575 5.495 1.955 ;
        RECT 4.905 1.065 5.075 1.395 ;
        RECT 5.325 1.035 5.495 1.575 ;
        RECT 5.665 1.385 5.835 2.135 ;
        RECT 6.005 2.105 6.175 2.375 ;
        RECT 6.410 2.355 6.740 2.635 ;
        RECT 6.995 2.105 7.165 2.375 ;
        RECT 7.375 2.175 7.745 2.635 ;
        RECT 6.005 1.935 7.165 2.105 ;
        RECT 7.970 2.005 8.140 2.465 ;
        RECT 8.320 2.125 9.190 2.465 ;
        RECT 9.360 2.195 9.610 2.635 ;
        RECT 9.015 2.115 9.190 2.125 ;
        RECT 9.015 2.035 9.210 2.115 ;
        RECT 7.455 1.835 8.140 2.005 ;
        RECT 8.310 1.935 8.840 1.955 ;
        RECT 7.455 1.765 7.715 1.835 ;
        RECT 6.285 1.595 7.715 1.765 ;
        RECT 8.310 1.665 8.870 1.935 ;
        RECT 5.665 1.215 7.375 1.385 ;
        RECT 4.565 0.715 5.145 0.895 ;
        RECT 2.915 0.255 3.850 0.425 ;
        RECT 4.445 0.085 4.775 0.540 ;
        RECT 4.975 0.505 5.145 0.715 ;
        RECT 5.325 0.705 5.975 1.035 ;
        RECT 4.975 0.335 5.315 0.505 ;
        RECT 6.165 0.475 6.335 1.215 ;
        RECT 6.505 0.765 7.035 1.045 ;
        RECT 7.205 1.005 7.375 1.215 ;
        RECT 7.545 0.835 7.715 1.595 ;
        RECT 5.485 0.305 6.335 0.475 ;
        RECT 6.915 0.085 7.245 0.545 ;
        RECT 7.455 0.445 7.715 0.835 ;
        RECT 7.885 1.655 8.870 1.665 ;
        RECT 9.040 1.745 9.210 2.035 ;
        RECT 9.780 2.085 9.950 2.375 ;
        RECT 10.120 2.255 10.450 2.635 ;
        RECT 9.780 1.915 10.545 2.085 ;
        RECT 7.885 1.495 8.520 1.655 ;
        RECT 9.040 1.575 10.205 1.745 ;
        RECT 7.885 0.705 8.095 1.495 ;
        RECT 9.040 1.485 9.210 1.575 ;
        RECT 8.405 0.920 8.575 1.325 ;
        RECT 8.745 1.315 9.210 1.485 ;
        RECT 10.375 1.325 10.545 1.915 ;
        RECT 10.720 1.495 10.970 2.635 ;
        RECT 8.745 0.535 8.915 1.315 ;
        RECT 10.375 1.295 11.020 1.325 ;
        RECT 9.125 0.865 9.295 1.145 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.125 0.695 9.655 0.865 ;
        RECT 7.455 0.275 7.785 0.445 ;
        RECT 8.005 0.255 8.915 0.535 ;
        RECT 9.085 0.085 9.255 0.525 ;
        RECT 9.485 0.465 9.655 0.695 ;
        RECT 9.825 0.635 10.115 1.065 ;
        RECT 10.345 0.995 11.020 1.295 ;
        RECT 10.345 0.465 10.515 0.995 ;
        RECT 9.485 0.295 10.515 0.465 ;
        RECT 10.720 0.085 10.890 0.545 ;
        RECT 0.000 -0.085 11.500 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 0.675 1.785 0.845 1.955 ;
        RECT 1.145 1.105 1.315 1.275 ;
        RECT 5.325 1.785 5.495 1.955 ;
        RECT 4.905 1.105 5.075 1.275 ;
        RECT 8.445 1.785 8.615 1.955 ;
        RECT 6.865 0.765 7.035 0.935 ;
        RECT 8.405 1.105 8.575 1.275 ;
        RECT 9.690 1.105 9.860 1.275 ;
        RECT 9.945 0.765 10.115 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
      LAYER met1 ;
        RECT 0.615 1.940 0.915 1.985 ;
        RECT 5.265 1.940 5.555 1.985 ;
        RECT 8.385 1.940 8.675 1.985 ;
        RECT 0.615 1.800 8.675 1.940 ;
        RECT 0.615 1.755 0.915 1.800 ;
        RECT 5.265 1.755 5.555 1.800 ;
        RECT 8.385 1.755 8.675 1.800 ;
        RECT 1.085 1.260 1.375 1.305 ;
        RECT 4.845 1.260 5.135 1.305 ;
        RECT 8.345 1.260 8.635 1.305 ;
        RECT 1.085 1.120 8.635 1.260 ;
        RECT 1.085 1.075 1.375 1.120 ;
        RECT 4.845 1.075 5.135 1.120 ;
        RECT 8.345 1.075 8.635 1.120 ;
  END
END sky130_fd_sc_hd__sdfrtn_1

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.500 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.975 0.490 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.144000 ;
    PORT
      LAYER li1 ;
        RECT 2.865 1.785 3.120 2.465 ;
        RECT 2.735 1.355 3.120 1.785 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 9.630 0.965 9.920 1.305 ;
        RECT 6.445 0.920 7.095 0.965 ;
        RECT 9.630 0.920 10.175 0.965 ;
        RECT 6.445 0.780 10.175 0.920 ;
        RECT 6.445 0.735 7.095 0.780 ;
        RECT 9.885 0.735 10.175 0.780 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.156600 ;
    PORT
      LAYER li1 ;
        RECT 4.020 0.710 4.395 1.700 ;
        RECT 4.020 0.285 4.275 0.710 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.730 2.465 ;
        RECT 1.485 1.070 1.730 1.985 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.500 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.880 1.355 1.015 ;
        RECT 2.305 0.880 3.640 1.145 ;
        RECT 0.005 0.725 4.885 0.880 ;
        RECT 6.955 0.785 7.865 1.005 ;
        RECT 10.550 0.785 11.480 1.015 ;
        RECT 5.935 0.725 11.480 0.785 ;
        RECT 0.005 0.465 11.480 0.725 ;
        RECT 0.005 0.200 2.295 0.465 ;
        RECT 3.150 0.200 11.480 0.465 ;
        RECT 0.005 0.105 1.355 0.200 ;
        RECT 4.895 0.105 11.480 0.200 ;
        RECT 0.215 -0.010 0.235 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.425 11.690 2.910 ;
        RECT -0.190 1.305 1.970 1.425 ;
        RECT 4.405 1.305 11.690 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.500 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 11.140 1.460 11.400 2.325 ;
        RECT 11.150 1.445 11.400 1.460 ;
        RECT 11.190 0.795 11.400 1.445 ;
        RECT 11.140 0.265 11.400 0.795 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.500 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.530 2.135 0.860 2.635 ;
        RECT 0.090 1.795 0.865 1.965 ;
        RECT 0.660 1.325 0.865 1.795 ;
        RECT 1.035 1.900 1.205 2.465 ;
        RECT 1.900 2.055 2.150 2.400 ;
        RECT 1.035 1.730 1.315 1.900 ;
        RECT 0.660 0.995 0.975 1.325 ;
        RECT 0.660 0.805 0.835 0.995 ;
        RECT 0.095 0.635 0.835 0.805 ;
        RECT 1.145 0.675 1.315 1.730 ;
        RECT 1.980 1.455 2.150 2.055 ;
        RECT 2.320 2.040 2.490 2.635 ;
        RECT 3.460 2.105 3.630 2.465 ;
        RECT 4.300 2.275 4.630 2.635 ;
        RECT 4.905 2.185 5.275 2.435 ;
        RECT 4.905 2.105 5.075 2.185 ;
        RECT 5.470 2.135 5.835 2.465 ;
        RECT 3.290 1.935 5.075 2.105 ;
        RECT 1.980 1.260 2.470 1.455 ;
        RECT 2.055 1.185 2.470 1.260 ;
        RECT 3.290 1.185 3.460 1.935 ;
        RECT 2.055 0.995 3.085 1.185 ;
        RECT 2.055 0.900 2.225 0.995 ;
        RECT 0.095 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.315 0.675 ;
        RECT 1.535 0.730 2.225 0.900 ;
        RECT 1.535 0.395 1.705 0.730 ;
        RECT 1.875 0.085 2.205 0.560 ;
        RECT 2.395 0.085 2.725 0.825 ;
        RECT 2.915 0.425 3.085 0.995 ;
        RECT 3.255 1.015 3.460 1.185 ;
        RECT 3.255 0.675 3.425 1.015 ;
        RECT 3.680 0.425 3.850 1.685 ;
        RECT 4.565 0.895 4.735 1.935 ;
        RECT 5.245 1.575 5.495 1.955 ;
        RECT 4.905 1.065 5.075 1.395 ;
        RECT 5.325 1.035 5.495 1.575 ;
        RECT 5.665 1.385 5.835 2.135 ;
        RECT 6.005 2.105 6.175 2.375 ;
        RECT 6.410 2.355 6.740 2.635 ;
        RECT 6.995 2.105 7.165 2.375 ;
        RECT 7.375 2.175 7.745 2.635 ;
        RECT 6.005 1.935 7.165 2.105 ;
        RECT 7.970 2.005 8.140 2.465 ;
        RECT 8.320 2.125 9.190 2.465 ;
        RECT 9.360 2.195 9.610 2.635 ;
        RECT 9.015 2.115 9.190 2.125 ;
        RECT 9.015 2.035 9.210 2.115 ;
        RECT 7.455 1.835 8.140 2.005 ;
        RECT 8.310 1.935 8.840 1.955 ;
        RECT 7.455 1.765 7.715 1.835 ;
        RECT 6.285 1.595 7.715 1.765 ;
        RECT 8.310 1.665 8.870 1.935 ;
        RECT 5.665 1.215 7.375 1.385 ;
        RECT 4.565 0.715 5.145 0.895 ;
        RECT 2.915 0.255 3.850 0.425 ;
        RECT 4.445 0.085 4.775 0.540 ;
        RECT 4.975 0.505 5.145 0.715 ;
        RECT 5.325 0.705 5.975 1.035 ;
        RECT 4.975 0.335 5.315 0.505 ;
        RECT 6.165 0.475 6.335 1.215 ;
        RECT 6.505 0.765 7.035 1.045 ;
        RECT 7.205 1.005 7.375 1.215 ;
        RECT 7.545 0.835 7.715 1.595 ;
        RECT 5.485 0.305 6.335 0.475 ;
        RECT 6.915 0.085 7.245 0.545 ;
        RECT 7.455 0.445 7.715 0.835 ;
        RECT 7.885 1.655 8.870 1.665 ;
        RECT 9.040 1.745 9.210 2.035 ;
        RECT 9.780 2.085 9.950 2.375 ;
        RECT 10.120 2.255 10.450 2.635 ;
        RECT 9.780 1.915 10.545 2.085 ;
        RECT 7.885 1.495 8.520 1.655 ;
        RECT 9.040 1.575 10.205 1.745 ;
        RECT 7.885 0.705 8.095 1.495 ;
        RECT 9.040 1.485 9.210 1.575 ;
        RECT 8.405 0.920 8.575 1.325 ;
        RECT 8.745 1.315 9.210 1.485 ;
        RECT 10.375 1.325 10.545 1.915 ;
        RECT 10.720 1.495 10.970 2.635 ;
        RECT 8.745 0.535 8.915 1.315 ;
        RECT 10.375 1.295 11.020 1.325 ;
        RECT 9.125 0.865 9.295 1.145 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.125 0.695 9.655 0.865 ;
        RECT 7.455 0.275 7.785 0.445 ;
        RECT 8.005 0.255 8.915 0.535 ;
        RECT 9.085 0.085 9.255 0.525 ;
        RECT 9.485 0.465 9.655 0.695 ;
        RECT 9.825 0.635 10.115 1.065 ;
        RECT 10.345 0.995 11.020 1.295 ;
        RECT 10.345 0.465 10.515 0.995 ;
        RECT 9.485 0.295 10.515 0.465 ;
        RECT 10.720 0.085 10.890 0.545 ;
        RECT 0.000 -0.085 11.500 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 1.035 1.785 1.205 1.955 ;
        RECT 0.805 1.105 0.975 1.275 ;
        RECT 5.325 1.785 5.495 1.955 ;
        RECT 4.905 1.105 5.075 1.275 ;
        RECT 8.445 1.785 8.615 1.955 ;
        RECT 6.865 0.765 7.035 0.935 ;
        RECT 8.405 1.105 8.575 1.275 ;
        RECT 9.690 1.105 9.860 1.275 ;
        RECT 9.945 0.765 10.115 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
      LAYER met1 ;
        RECT 0.970 1.940 1.270 1.985 ;
        RECT 5.265 1.940 5.555 1.985 ;
        RECT 8.385 1.940 8.675 1.985 ;
        RECT 0.970 1.800 8.675 1.940 ;
        RECT 0.970 1.755 1.270 1.800 ;
        RECT 5.265 1.755 5.555 1.800 ;
        RECT 8.385 1.755 8.675 1.800 ;
        RECT 0.745 1.260 1.035 1.305 ;
        RECT 4.845 1.260 5.135 1.305 ;
        RECT 8.345 1.260 8.635 1.305 ;
        RECT 0.745 1.120 8.635 1.260 ;
        RECT 0.745 1.075 1.035 1.120 ;
        RECT 4.845 1.075 5.135 1.120 ;
        RECT 8.345 1.075 8.635 1.120 ;
  END
END sky130_fd_sc_hd__sdfrtp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfrtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.960 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.975 0.490 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.144000 ;
    PORT
      LAYER li1 ;
        RECT 2.865 1.785 3.120 2.465 ;
        RECT 2.735 1.355 3.120 1.785 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 9.630 0.965 9.920 1.305 ;
        RECT 6.445 0.920 7.095 0.965 ;
        RECT 9.630 0.920 10.175 0.965 ;
        RECT 6.445 0.780 10.175 0.920 ;
        RECT 6.445 0.735 7.095 0.780 ;
        RECT 9.885 0.735 10.175 0.780 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.156600 ;
    PORT
      LAYER li1 ;
        RECT 4.020 0.710 4.395 1.700 ;
        RECT 4.020 0.285 4.275 0.710 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.730 2.465 ;
        RECT 1.485 1.070 1.730 1.985 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.960 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.880 1.355 1.015 ;
        RECT 2.305 0.880 3.640 1.145 ;
        RECT 0.005 0.725 4.885 0.880 ;
        RECT 6.955 0.785 7.865 1.005 ;
        RECT 10.550 0.785 11.910 1.015 ;
        RECT 5.935 0.725 11.910 0.785 ;
        RECT 0.005 0.465 11.910 0.725 ;
        RECT 0.005 0.200 2.295 0.465 ;
        RECT 3.150 0.200 11.910 0.465 ;
        RECT 0.005 0.105 1.355 0.200 ;
        RECT 4.895 0.105 11.910 0.200 ;
        RECT 0.215 -0.010 0.235 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.425 12.150 2.910 ;
        RECT -0.190 1.305 1.970 1.425 ;
        RECT 4.405 1.305 12.150 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.960 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 11.140 1.460 11.400 2.325 ;
        RECT 11.150 1.445 11.400 1.460 ;
        RECT 11.190 0.795 11.400 1.445 ;
        RECT 11.140 0.265 11.400 0.795 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.960 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.530 2.135 0.860 2.635 ;
        RECT 0.090 1.795 0.865 1.965 ;
        RECT 0.660 1.325 0.865 1.795 ;
        RECT 1.035 1.900 1.205 2.465 ;
        RECT 1.900 2.055 2.150 2.400 ;
        RECT 1.035 1.730 1.315 1.900 ;
        RECT 0.660 0.995 0.975 1.325 ;
        RECT 0.660 0.805 0.835 0.995 ;
        RECT 0.095 0.635 0.835 0.805 ;
        RECT 1.145 0.675 1.315 1.730 ;
        RECT 1.980 1.455 2.150 2.055 ;
        RECT 2.320 2.040 2.490 2.635 ;
        RECT 3.460 2.105 3.630 2.465 ;
        RECT 4.300 2.275 4.630 2.635 ;
        RECT 4.905 2.185 5.275 2.435 ;
        RECT 4.905 2.105 5.075 2.185 ;
        RECT 5.470 2.135 5.835 2.465 ;
        RECT 3.290 1.935 5.075 2.105 ;
        RECT 1.980 1.260 2.470 1.455 ;
        RECT 2.055 1.185 2.470 1.260 ;
        RECT 3.290 1.185 3.460 1.935 ;
        RECT 2.055 0.995 3.085 1.185 ;
        RECT 2.055 0.900 2.225 0.995 ;
        RECT 0.095 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.315 0.675 ;
        RECT 1.535 0.730 2.225 0.900 ;
        RECT 1.535 0.395 1.705 0.730 ;
        RECT 1.875 0.085 2.205 0.560 ;
        RECT 2.395 0.085 2.725 0.825 ;
        RECT 2.915 0.425 3.085 0.995 ;
        RECT 3.255 1.015 3.460 1.185 ;
        RECT 3.255 0.675 3.425 1.015 ;
        RECT 3.680 0.425 3.850 1.685 ;
        RECT 4.565 0.895 4.735 1.935 ;
        RECT 5.245 1.575 5.495 1.955 ;
        RECT 4.905 1.065 5.075 1.395 ;
        RECT 5.325 1.035 5.495 1.575 ;
        RECT 5.665 1.385 5.835 2.135 ;
        RECT 6.005 2.105 6.175 2.375 ;
        RECT 6.410 2.355 6.740 2.635 ;
        RECT 6.995 2.105 7.165 2.375 ;
        RECT 7.375 2.175 7.745 2.635 ;
        RECT 6.005 1.935 7.165 2.105 ;
        RECT 7.970 2.005 8.140 2.465 ;
        RECT 8.320 2.125 9.190 2.465 ;
        RECT 9.360 2.195 9.610 2.635 ;
        RECT 9.015 2.115 9.190 2.125 ;
        RECT 9.015 2.035 9.210 2.115 ;
        RECT 7.455 1.835 8.140 2.005 ;
        RECT 8.310 1.935 8.840 1.955 ;
        RECT 7.455 1.765 7.715 1.835 ;
        RECT 6.285 1.595 7.715 1.765 ;
        RECT 8.310 1.665 8.870 1.935 ;
        RECT 5.665 1.215 7.375 1.385 ;
        RECT 4.565 0.715 5.145 0.895 ;
        RECT 2.915 0.255 3.850 0.425 ;
        RECT 4.445 0.085 4.775 0.540 ;
        RECT 4.975 0.505 5.145 0.715 ;
        RECT 5.325 0.705 5.975 1.035 ;
        RECT 4.975 0.335 5.315 0.505 ;
        RECT 6.165 0.475 6.335 1.215 ;
        RECT 6.505 0.765 7.035 1.045 ;
        RECT 7.205 1.005 7.375 1.215 ;
        RECT 7.545 0.835 7.715 1.595 ;
        RECT 5.485 0.305 6.335 0.475 ;
        RECT 6.915 0.085 7.245 0.545 ;
        RECT 7.455 0.445 7.715 0.835 ;
        RECT 7.885 1.655 8.870 1.665 ;
        RECT 9.040 1.745 9.210 2.035 ;
        RECT 9.780 2.085 9.950 2.375 ;
        RECT 10.120 2.255 10.450 2.635 ;
        RECT 9.780 1.915 10.545 2.085 ;
        RECT 7.885 1.495 8.520 1.655 ;
        RECT 9.040 1.575 10.205 1.745 ;
        RECT 7.885 0.705 8.095 1.495 ;
        RECT 9.040 1.485 9.210 1.575 ;
        RECT 8.405 0.920 8.575 1.325 ;
        RECT 8.745 1.315 9.210 1.485 ;
        RECT 10.375 1.325 10.545 1.915 ;
        RECT 10.720 1.495 10.970 2.635 ;
        RECT 11.570 1.495 11.820 2.635 ;
        RECT 8.745 0.535 8.915 1.315 ;
        RECT 10.375 1.295 11.020 1.325 ;
        RECT 9.125 0.865 9.295 1.145 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.125 0.695 9.655 0.865 ;
        RECT 7.455 0.275 7.785 0.445 ;
        RECT 8.005 0.255 8.915 0.535 ;
        RECT 9.085 0.085 9.255 0.525 ;
        RECT 9.485 0.465 9.655 0.695 ;
        RECT 9.825 0.635 10.115 1.065 ;
        RECT 10.345 0.995 11.020 1.295 ;
        RECT 10.345 0.465 10.515 0.995 ;
        RECT 9.485 0.295 10.515 0.465 ;
        RECT 10.720 0.085 10.890 0.545 ;
        RECT 11.570 0.085 11.740 0.545 ;
        RECT 0.000 -0.085 11.960 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 1.035 1.785 1.205 1.955 ;
        RECT 0.805 1.105 0.975 1.275 ;
        RECT 5.325 1.785 5.495 1.955 ;
        RECT 4.905 1.105 5.075 1.275 ;
        RECT 8.445 1.785 8.615 1.955 ;
        RECT 6.865 0.765 7.035 0.935 ;
        RECT 8.405 1.105 8.575 1.275 ;
        RECT 9.690 1.105 9.860 1.275 ;
        RECT 9.945 0.765 10.115 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
      LAYER met1 ;
        RECT 0.970 1.940 1.270 1.985 ;
        RECT 5.265 1.940 5.555 1.985 ;
        RECT 8.385 1.940 8.675 1.985 ;
        RECT 0.970 1.800 8.675 1.940 ;
        RECT 0.970 1.755 1.270 1.800 ;
        RECT 5.265 1.755 5.555 1.800 ;
        RECT 8.385 1.755 8.675 1.800 ;
        RECT 0.745 1.260 1.035 1.305 ;
        RECT 4.845 1.260 5.135 1.305 ;
        RECT 8.345 1.260 8.635 1.305 ;
        RECT 0.745 1.120 8.635 1.260 ;
        RECT 0.745 1.075 1.035 1.120 ;
        RECT 4.845 1.075 5.135 1.120 ;
        RECT 8.345 1.075 8.635 1.120 ;
  END
END sky130_fd_sc_hd__sdfrtp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfrtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER li1 ;
        RECT 0.140 0.975 0.490 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.144000 ;
    PORT
      LAYER li1 ;
        RECT 2.865 1.785 3.120 2.465 ;
        RECT 2.735 1.355 3.120 1.785 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 9.630 0.965 9.920 1.305 ;
        RECT 6.445 0.920 7.095 0.965 ;
        RECT 9.630 0.920 10.175 0.965 ;
        RECT 6.445 0.780 10.175 0.920 ;
        RECT 6.445 0.735 7.095 0.780 ;
        RECT 9.885 0.735 10.175 0.780 ;
    END
  END RESET_B
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.156600 ;
    PORT
      LAYER li1 ;
        RECT 4.020 0.710 4.395 1.700 ;
        RECT 4.020 0.285 4.275 0.710 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.435000 ;
    PORT
      LAYER li1 ;
        RECT 1.465 1.985 1.730 2.465 ;
        RECT 1.485 1.070 1.730 1.985 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.880 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.880 1.355 1.015 ;
        RECT 2.305 0.880 3.640 1.145 ;
        RECT 0.005 0.725 4.885 0.880 ;
        RECT 6.955 0.785 7.865 1.005 ;
        RECT 10.550 0.785 12.750 1.015 ;
        RECT 5.935 0.725 12.750 0.785 ;
        RECT 0.005 0.465 12.750 0.725 ;
        RECT 0.005 0.200 2.295 0.465 ;
        RECT 3.150 0.200 12.750 0.465 ;
        RECT 0.005 0.105 1.355 0.200 ;
        RECT 4.895 0.105 12.750 0.200 ;
        RECT 0.215 -0.010 0.235 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.425 13.070 2.910 ;
        RECT -0.190 1.305 1.970 1.425 ;
        RECT 4.405 1.305 13.070 1.425 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 12.880 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 11.140 1.460 11.400 2.325 ;
        RECT 11.150 1.445 11.400 1.460 ;
        RECT 11.190 1.325 11.400 1.445 ;
        RECT 11.990 1.325 12.240 2.325 ;
        RECT 11.190 0.995 12.240 1.325 ;
        RECT 11.190 0.795 11.400 0.995 ;
        RECT 11.140 0.265 11.400 0.795 ;
        RECT 11.990 0.265 12.240 0.995 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 12.880 2.805 ;
        RECT 0.090 1.965 0.345 2.465 ;
        RECT 0.530 2.135 0.860 2.635 ;
        RECT 0.090 1.795 0.865 1.965 ;
        RECT 0.660 1.325 0.865 1.795 ;
        RECT 1.035 1.900 1.205 2.465 ;
        RECT 1.900 2.055 2.150 2.400 ;
        RECT 1.035 1.730 1.315 1.900 ;
        RECT 0.660 0.995 0.975 1.325 ;
        RECT 0.660 0.805 0.835 0.995 ;
        RECT 0.095 0.635 0.835 0.805 ;
        RECT 1.145 0.675 1.315 1.730 ;
        RECT 1.980 1.455 2.150 2.055 ;
        RECT 2.320 2.040 2.490 2.635 ;
        RECT 3.460 2.105 3.630 2.465 ;
        RECT 4.300 2.275 4.630 2.635 ;
        RECT 4.905 2.185 5.275 2.435 ;
        RECT 4.905 2.105 5.075 2.185 ;
        RECT 5.470 2.135 5.835 2.465 ;
        RECT 3.290 1.935 5.075 2.105 ;
        RECT 1.980 1.260 2.470 1.455 ;
        RECT 2.055 1.185 2.470 1.260 ;
        RECT 3.290 1.185 3.460 1.935 ;
        RECT 2.055 0.995 3.085 1.185 ;
        RECT 2.055 0.900 2.225 0.995 ;
        RECT 0.095 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.315 0.675 ;
        RECT 1.535 0.730 2.225 0.900 ;
        RECT 1.535 0.395 1.705 0.730 ;
        RECT 1.875 0.085 2.205 0.560 ;
        RECT 2.395 0.085 2.725 0.825 ;
        RECT 2.915 0.425 3.085 0.995 ;
        RECT 3.255 1.015 3.460 1.185 ;
        RECT 3.255 0.675 3.425 1.015 ;
        RECT 3.680 0.425 3.850 1.685 ;
        RECT 4.565 0.895 4.735 1.935 ;
        RECT 5.245 1.575 5.495 1.955 ;
        RECT 4.905 1.065 5.075 1.395 ;
        RECT 5.325 1.035 5.495 1.575 ;
        RECT 5.665 1.385 5.835 2.135 ;
        RECT 6.005 2.105 6.175 2.375 ;
        RECT 6.410 2.355 6.740 2.635 ;
        RECT 6.995 2.105 7.165 2.375 ;
        RECT 7.375 2.175 7.745 2.635 ;
        RECT 6.005 1.935 7.165 2.105 ;
        RECT 7.970 2.005 8.140 2.465 ;
        RECT 8.320 2.125 9.190 2.465 ;
        RECT 9.360 2.195 9.610 2.635 ;
        RECT 9.015 2.115 9.190 2.125 ;
        RECT 9.015 2.035 9.210 2.115 ;
        RECT 7.455 1.835 8.140 2.005 ;
        RECT 8.310 1.935 8.840 1.955 ;
        RECT 7.455 1.765 7.715 1.835 ;
        RECT 6.285 1.595 7.715 1.765 ;
        RECT 8.310 1.665 8.870 1.935 ;
        RECT 5.665 1.215 7.375 1.385 ;
        RECT 4.565 0.715 5.145 0.895 ;
        RECT 2.915 0.255 3.850 0.425 ;
        RECT 4.445 0.085 4.775 0.540 ;
        RECT 4.975 0.505 5.145 0.715 ;
        RECT 5.325 0.705 5.975 1.035 ;
        RECT 4.975 0.335 5.315 0.505 ;
        RECT 6.165 0.475 6.335 1.215 ;
        RECT 6.505 0.765 7.035 1.045 ;
        RECT 7.205 1.005 7.375 1.215 ;
        RECT 7.545 0.835 7.715 1.595 ;
        RECT 5.485 0.305 6.335 0.475 ;
        RECT 6.915 0.085 7.245 0.545 ;
        RECT 7.455 0.445 7.715 0.835 ;
        RECT 7.885 1.655 8.870 1.665 ;
        RECT 9.040 1.745 9.210 2.035 ;
        RECT 9.780 2.085 9.950 2.375 ;
        RECT 10.120 2.255 10.450 2.635 ;
        RECT 9.780 1.915 10.545 2.085 ;
        RECT 7.885 1.495 8.520 1.655 ;
        RECT 9.040 1.575 10.205 1.745 ;
        RECT 7.885 0.705 8.095 1.495 ;
        RECT 9.040 1.485 9.210 1.575 ;
        RECT 8.405 0.920 8.575 1.325 ;
        RECT 8.745 1.315 9.210 1.485 ;
        RECT 10.375 1.325 10.545 1.915 ;
        RECT 10.720 1.495 10.970 2.635 ;
        RECT 11.570 1.495 11.820 2.635 ;
        RECT 12.410 1.495 12.660 2.635 ;
        RECT 8.745 0.535 8.915 1.315 ;
        RECT 10.375 1.295 11.020 1.325 ;
        RECT 9.125 0.865 9.295 1.145 ;
        RECT 9.525 1.065 10.115 1.275 ;
        RECT 9.125 0.695 9.655 0.865 ;
        RECT 7.455 0.275 7.785 0.445 ;
        RECT 8.005 0.255 8.915 0.535 ;
        RECT 9.085 0.085 9.255 0.525 ;
        RECT 9.485 0.465 9.655 0.695 ;
        RECT 9.825 0.635 10.115 1.065 ;
        RECT 10.345 0.995 11.020 1.295 ;
        RECT 10.345 0.465 10.515 0.995 ;
        RECT 9.485 0.295 10.515 0.465 ;
        RECT 10.720 0.085 10.890 0.545 ;
        RECT 11.570 0.085 11.740 0.545 ;
        RECT 12.410 0.085 12.580 0.545 ;
        RECT 0.000 -0.085 12.880 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 1.035 1.785 1.205 1.955 ;
        RECT 0.805 1.105 0.975 1.275 ;
        RECT 5.325 1.785 5.495 1.955 ;
        RECT 4.905 1.105 5.075 1.275 ;
        RECT 8.445 1.785 8.615 1.955 ;
        RECT 6.865 0.765 7.035 0.935 ;
        RECT 8.405 1.105 8.575 1.275 ;
        RECT 9.690 1.105 9.860 1.275 ;
        RECT 9.945 0.765 10.115 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
      LAYER met1 ;
        RECT 0.970 1.940 1.270 1.985 ;
        RECT 5.265 1.940 5.555 1.985 ;
        RECT 8.385 1.940 8.675 1.985 ;
        RECT 0.970 1.800 8.675 1.940 ;
        RECT 0.970 1.755 1.270 1.800 ;
        RECT 5.265 1.755 5.555 1.800 ;
        RECT 8.385 1.755 8.675 1.800 ;
        RECT 0.745 1.260 1.035 1.305 ;
        RECT 4.845 1.260 5.135 1.305 ;
        RECT 8.345 1.260 8.635 1.305 ;
        RECT 0.745 1.120 8.635 1.260 ;
        RECT 0.745 1.075 1.035 1.120 ;
        RECT 4.845 1.075 5.135 1.120 ;
        RECT 8.345 1.075 8.635 1.120 ;
  END
END sky130_fd_sc_hd__sdfrtp_4

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfsbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.340 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.590 3.085 1.960 ;
        RECT 2.905 1.055 3.565 1.590 ;
        RECT 2.905 0.725 3.100 1.055 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.055 0.765 1.335 1.675 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.345 1.675 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER met1 ;
        RECT 0.550 1.260 0.840 1.305 ;
        RECT 2.385 1.260 2.675 1.305 ;
        RECT 0.550 1.120 2.675 1.260 ;
        RECT 0.550 1.075 0.840 1.120 ;
        RECT 2.385 1.075 2.675 1.120 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 6.580 1.600 6.870 1.645 ;
        RECT 8.825 1.600 9.115 1.645 ;
        RECT 6.580 1.460 9.115 1.600 ;
        RECT 6.580 1.415 6.870 1.460 ;
        RECT 8.825 1.415 9.115 1.460 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 13.340 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 7.040 0.785 8.795 1.005 ;
        RECT 10.990 0.785 13.335 1.015 ;
        RECT 0.005 0.105 13.335 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 13.530 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 13.340 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 12.915 1.495 13.255 2.450 ;
        RECT 13.070 0.825 13.255 1.495 ;
        RECT 12.915 0.275 13.255 0.825 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 11.500 0.255 11.830 2.465 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 13.340 2.805 ;
        RECT 0.085 2.025 0.345 2.465 ;
        RECT 0.515 2.195 0.765 2.635 ;
        RECT 0.935 2.255 2.045 2.465 ;
        RECT 0.935 2.025 1.105 2.255 ;
        RECT 2.270 2.085 2.520 2.465 ;
        RECT 2.690 2.140 3.030 2.635 ;
        RECT 0.085 1.845 1.105 2.025 ;
        RECT 1.295 1.870 1.695 2.075 ;
        RECT 0.545 0.765 0.825 1.675 ;
        RECT 1.505 0.705 1.695 1.870 ;
        RECT 1.865 1.770 2.520 2.085 ;
        RECT 3.255 1.955 3.425 2.325 ;
        RECT 3.595 2.275 3.925 2.635 ;
        RECT 4.095 2.135 4.440 2.465 ;
        RECT 3.255 1.775 3.995 1.955 ;
        RECT 1.865 0.905 2.200 1.770 ;
        RECT 2.370 1.075 2.700 1.600 ;
        RECT 1.865 0.715 2.515 0.905 ;
        RECT 3.735 0.885 3.995 1.775 ;
        RECT 1.495 0.665 1.695 0.705 ;
        RECT 1.475 0.655 1.695 0.665 ;
        RECT 1.475 0.645 1.670 0.655 ;
        RECT 1.460 0.635 1.670 0.645 ;
        RECT 1.445 0.630 1.670 0.635 ;
        RECT 1.440 0.620 1.670 0.630 ;
        RECT 1.430 0.615 1.670 0.620 ;
        RECT 1.420 0.610 1.660 0.615 ;
        RECT 1.405 0.605 1.660 0.610 ;
        RECT 1.395 0.600 1.660 0.605 ;
        RECT 0.085 0.085 0.480 0.595 ;
        RECT 1.380 0.590 1.660 0.600 ;
        RECT 1.380 0.560 1.655 0.590 ;
        RECT 0.875 0.280 1.655 0.560 ;
        RECT 1.825 0.085 2.005 0.545 ;
        RECT 2.260 0.255 2.515 0.715 ;
        RECT 3.270 0.715 3.995 0.885 ;
        RECT 4.165 1.420 4.440 2.135 ;
        RECT 4.610 1.615 4.830 2.465 ;
        RECT 5.030 2.135 5.755 2.465 ;
        RECT 5.945 2.275 6.275 2.635 ;
        RECT 4.610 1.590 4.915 1.615 ;
        RECT 4.660 1.445 4.915 1.590 ;
        RECT 5.205 1.575 5.415 1.955 ;
        RECT 4.165 1.090 4.490 1.420 ;
        RECT 2.690 0.085 3.030 0.555 ;
        RECT 3.270 0.255 3.455 0.715 ;
        RECT 4.165 0.585 4.335 1.090 ;
        RECT 4.660 0.920 4.830 1.445 ;
        RECT 5.585 1.395 5.755 2.135 ;
        RECT 6.550 2.105 6.765 2.450 ;
        RECT 7.005 2.125 7.960 2.635 ;
        RECT 8.130 2.125 8.935 2.460 ;
        RECT 9.195 2.235 9.525 2.635 ;
        RECT 5.925 1.935 6.765 2.105 ;
        RECT 8.765 2.065 8.935 2.125 ;
        RECT 9.695 2.065 9.910 2.450 ;
        RECT 10.135 2.235 10.465 2.635 ;
        RECT 5.925 1.575 6.095 1.935 ;
        RECT 6.640 1.445 7.015 1.765 ;
        RECT 7.190 1.495 8.005 1.955 ;
        RECT 5.085 1.275 6.435 1.395 ;
        RECT 7.300 1.275 7.660 1.325 ;
        RECT 3.630 0.085 3.940 0.545 ;
        RECT 4.110 0.255 4.335 0.585 ;
        RECT 4.505 0.255 4.830 0.920 ;
        RECT 5.000 1.225 7.660 1.275 ;
        RECT 5.000 0.255 5.440 1.225 ;
        RECT 5.610 0.805 5.975 1.015 ;
        RECT 6.250 0.975 7.660 1.225 ;
        RECT 7.835 0.895 8.005 1.495 ;
        RECT 8.365 1.075 8.595 1.905 ;
        RECT 8.765 1.895 10.465 2.065 ;
        RECT 8.885 1.525 10.075 1.725 ;
        RECT 10.245 1.525 10.465 1.895 ;
        RECT 8.885 1.415 9.110 1.525 ;
        RECT 10.635 1.355 10.895 2.465 ;
        RECT 11.120 1.485 11.330 2.635 ;
        RECT 8.810 0.895 9.040 1.245 ;
        RECT 5.610 0.635 6.535 0.805 ;
        RECT 5.610 0.085 6.095 0.465 ;
        RECT 6.275 0.255 6.535 0.635 ;
        RECT 6.735 0.085 7.630 0.805 ;
        RECT 7.835 0.695 9.040 0.895 ;
        RECT 9.290 1.185 10.895 1.355 ;
        RECT 9.290 0.855 9.465 1.185 ;
        RECT 9.655 0.845 10.545 1.015 ;
        RECT 9.655 0.445 9.825 0.845 ;
        RECT 8.410 0.275 9.825 0.445 ;
        RECT 10.220 0.085 10.390 0.545 ;
        RECT 10.715 0.540 10.895 1.185 ;
        RECT 12.060 1.325 12.270 2.465 ;
        RECT 12.575 1.575 12.745 2.635 ;
        RECT 12.060 0.995 12.900 1.325 ;
        RECT 10.560 0.255 10.895 0.540 ;
        RECT 11.120 0.085 11.330 0.885 ;
        RECT 12.060 0.255 12.270 0.995 ;
        RECT 12.540 0.085 12.745 0.825 ;
        RECT 0.000 -0.085 13.340 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 0.610 1.105 0.780 1.275 ;
        RECT 1.525 1.445 1.695 1.615 ;
        RECT 3.825 1.785 3.995 1.955 ;
        RECT 2.445 1.105 2.615 1.275 ;
        RECT 5.205 1.785 5.375 1.955 ;
        RECT 4.745 1.445 4.915 1.615 ;
        RECT 4.285 1.105 4.455 1.275 ;
        RECT 7.505 1.785 7.675 1.955 ;
        RECT 8.885 1.445 9.055 1.615 ;
        RECT 8.425 1.105 8.595 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
      LAYER met1 ;
        RECT 3.765 1.940 4.055 1.985 ;
        RECT 5.145 1.940 5.435 1.985 ;
        RECT 7.445 1.940 7.735 1.985 ;
        RECT 3.765 1.800 7.735 1.940 ;
        RECT 3.765 1.755 4.055 1.800 ;
        RECT 5.145 1.755 5.435 1.800 ;
        RECT 7.445 1.755 7.735 1.800 ;
        RECT 1.465 1.600 1.755 1.645 ;
        RECT 4.685 1.600 4.975 1.645 ;
        RECT 1.465 1.460 4.975 1.600 ;
        RECT 1.465 1.415 1.755 1.460 ;
        RECT 4.685 1.415 4.975 1.460 ;
        RECT 4.225 1.260 4.515 1.305 ;
        RECT 8.365 1.260 8.655 1.305 ;
        RECT 4.225 1.120 8.655 1.260 ;
        RECT 4.225 1.075 4.515 1.120 ;
        RECT 8.365 1.075 8.655 1.120 ;
  END
END sky130_fd_sc_hd__sdfsbp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfsbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfsbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.260 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.615 3.100 1.970 ;
        RECT 2.905 1.055 3.565 1.615 ;
        RECT 2.905 0.725 3.100 1.055 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.050 0.765 1.335 1.675 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.340 1.675 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER met1 ;
        RECT 0.545 1.260 0.835 1.305 ;
        RECT 2.385 1.260 2.675 1.305 ;
        RECT 0.545 1.120 2.675 1.260 ;
        RECT 0.545 1.075 0.835 1.120 ;
        RECT 2.385 1.075 2.675 1.120 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 6.580 1.600 6.870 1.645 ;
        RECT 8.880 1.600 9.170 1.645 ;
        RECT 6.580 1.460 9.170 1.600 ;
        RECT 6.580 1.415 6.870 1.460 ;
        RECT 8.880 1.415 9.170 1.460 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 14.260 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 7.055 0.785 8.845 1.005 ;
        RECT 10.950 0.785 14.250 1.015 ;
        RECT 0.005 0.105 14.250 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 14.450 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 14.260 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 13.410 1.495 13.740 2.450 ;
        RECT 13.515 0.825 13.740 1.495 ;
        RECT 13.410 0.275 13.740 0.825 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 11.460 0.255 11.855 2.465 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 14.260 2.805 ;
        RECT 0.085 2.075 0.345 2.465 ;
        RECT 0.515 2.275 0.845 2.635 ;
        RECT 1.015 2.255 2.105 2.465 ;
        RECT 1.015 2.075 1.185 2.255 ;
        RECT 2.275 2.085 2.535 2.465 ;
        RECT 2.705 2.140 3.100 2.635 ;
        RECT 0.085 1.845 1.185 2.075 ;
        RECT 1.355 1.845 1.695 2.085 ;
        RECT 0.540 0.765 0.820 1.675 ;
        RECT 1.505 0.720 1.695 1.845 ;
        RECT 1.500 0.705 1.695 0.720 ;
        RECT 1.980 1.760 2.535 2.085 ;
        RECT 3.270 2.000 3.475 2.325 ;
        RECT 3.645 2.275 3.975 2.635 ;
        RECT 4.145 2.135 4.440 2.465 ;
        RECT 3.270 1.830 3.995 2.000 ;
        RECT 1.980 0.905 2.235 1.760 ;
        RECT 2.405 1.075 2.735 1.590 ;
        RECT 1.980 0.715 2.530 0.905 ;
        RECT 3.735 0.885 3.995 1.830 ;
        RECT 1.495 0.645 1.695 0.705 ;
        RECT 1.495 0.595 1.670 0.645 ;
        RECT 0.085 0.085 0.700 0.595 ;
        RECT 0.870 0.255 1.670 0.595 ;
        RECT 1.840 0.085 2.090 0.545 ;
        RECT 2.260 0.255 2.530 0.715 ;
        RECT 3.270 0.715 3.995 0.885 ;
        RECT 4.165 1.420 4.440 2.135 ;
        RECT 4.665 1.615 4.890 2.465 ;
        RECT 5.060 2.135 5.805 2.465 ;
        RECT 6.000 2.275 6.330 2.635 ;
        RECT 4.665 1.590 4.970 1.615 ;
        RECT 4.715 1.445 4.970 1.590 ;
        RECT 5.205 1.575 5.465 1.955 ;
        RECT 4.165 1.090 4.490 1.420 ;
        RECT 2.700 0.085 3.100 0.555 ;
        RECT 3.270 0.255 3.470 0.715 ;
        RECT 4.165 0.585 4.335 1.090 ;
        RECT 4.715 0.920 4.885 1.445 ;
        RECT 5.635 1.395 5.805 2.135 ;
        RECT 6.605 2.105 6.820 2.450 ;
        RECT 7.060 2.125 8.015 2.635 ;
        RECT 8.185 2.125 8.990 2.460 ;
        RECT 9.160 2.235 9.490 2.635 ;
        RECT 5.975 1.935 6.820 2.105 ;
        RECT 8.820 2.065 8.990 2.125 ;
        RECT 9.660 2.065 9.930 2.450 ;
        RECT 10.100 2.235 10.430 2.635 ;
        RECT 5.975 1.575 6.145 1.935 ;
        RECT 6.640 1.445 7.065 1.765 ;
        RECT 7.385 1.705 8.055 1.955 ;
        RECT 5.140 1.275 6.475 1.395 ;
        RECT 7.355 1.275 7.705 1.325 ;
        RECT 3.640 0.085 3.940 0.545 ;
        RECT 4.110 0.255 4.335 0.585 ;
        RECT 4.505 0.255 4.885 0.920 ;
        RECT 5.055 1.225 7.705 1.275 ;
        RECT 5.055 0.255 5.450 1.225 ;
        RECT 5.620 0.805 6.015 1.015 ;
        RECT 6.305 0.975 7.705 1.225 ;
        RECT 7.885 0.895 8.055 1.705 ;
        RECT 8.420 1.075 8.650 1.905 ;
        RECT 8.820 1.895 10.430 2.065 ;
        RECT 8.880 1.525 9.935 1.725 ;
        RECT 10.105 1.525 10.430 1.895 ;
        RECT 8.880 1.435 9.115 1.525 ;
        RECT 10.600 1.355 10.845 2.465 ;
        RECT 11.080 1.485 11.290 2.635 ;
        RECT 12.025 1.485 12.315 2.635 ;
        RECT 8.830 0.895 9.085 1.265 ;
        RECT 5.620 0.635 6.550 0.805 ;
        RECT 5.665 0.085 6.165 0.465 ;
        RECT 6.335 0.255 6.550 0.635 ;
        RECT 6.720 0.085 7.705 0.805 ;
        RECT 7.885 0.695 9.085 0.895 ;
        RECT 9.285 1.185 10.910 1.355 ;
        RECT 9.285 0.855 9.515 1.185 ;
        RECT 9.685 0.845 10.560 1.015 ;
        RECT 9.685 0.515 9.855 0.845 ;
        RECT 10.730 0.585 10.910 1.185 ;
        RECT 12.530 1.325 12.715 2.465 ;
        RECT 12.885 1.635 13.240 2.635 ;
        RECT 13.910 1.485 14.175 2.635 ;
        RECT 12.530 0.995 13.345 1.325 ;
        RECT 8.465 0.275 9.855 0.515 ;
        RECT 10.035 0.085 10.285 0.545 ;
        RECT 10.465 0.255 10.910 0.585 ;
        RECT 11.120 0.085 11.290 0.885 ;
        RECT 12.025 0.085 12.315 0.885 ;
        RECT 12.530 0.255 12.715 0.995 ;
        RECT 12.885 0.085 13.240 0.825 ;
        RECT 13.910 0.085 14.175 0.885 ;
        RECT 0.000 -0.085 14.260 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 0.605 1.105 0.775 1.275 ;
        RECT 1.525 1.445 1.695 1.615 ;
        RECT 3.825 1.785 3.995 1.955 ;
        RECT 2.445 1.105 2.615 1.275 ;
        RECT 5.260 1.785 5.430 1.955 ;
        RECT 4.800 1.445 4.970 1.615 ;
        RECT 4.285 1.105 4.455 1.275 ;
        RECT 7.560 1.785 7.730 1.955 ;
        RECT 8.940 1.445 9.110 1.615 ;
        RECT 8.480 1.105 8.650 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
      LAYER met1 ;
        RECT 3.765 1.940 4.055 1.985 ;
        RECT 5.200 1.940 5.490 1.985 ;
        RECT 7.500 1.940 7.790 1.985 ;
        RECT 3.765 1.800 7.790 1.940 ;
        RECT 3.765 1.755 4.055 1.800 ;
        RECT 5.200 1.755 5.490 1.800 ;
        RECT 7.500 1.755 7.790 1.800 ;
        RECT 1.465 1.600 1.755 1.645 ;
        RECT 4.740 1.600 5.030 1.645 ;
        RECT 1.465 1.460 5.030 1.600 ;
        RECT 1.465 1.415 1.755 1.460 ;
        RECT 4.740 1.415 5.030 1.460 ;
        RECT 4.225 1.260 4.515 1.305 ;
        RECT 8.420 1.260 8.710 1.305 ;
        RECT 4.225 1.120 8.710 1.260 ;
        RECT 4.225 1.075 4.515 1.120 ;
        RECT 8.420 1.075 8.710 1.120 ;
  END
END sky130_fd_sc_hd__sdfsbp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfstp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.420 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.615 3.085 1.960 ;
        RECT 2.905 1.055 3.565 1.615 ;
        RECT 2.905 0.725 3.100 1.055 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.050 0.765 1.335 1.675 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.340 1.675 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER met1 ;
        RECT 0.545 1.260 0.835 1.305 ;
        RECT 2.385 1.260 2.675 1.305 ;
        RECT 0.545 1.120 2.675 1.260 ;
        RECT 0.545 1.075 0.835 1.120 ;
        RECT 2.385 1.075 2.675 1.120 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 6.580 1.600 6.870 1.645 ;
        RECT 8.880 1.600 9.170 1.645 ;
        RECT 6.580 1.460 9.170 1.600 ;
        RECT 6.580 1.415 6.870 1.460 ;
        RECT 8.880 1.415 9.170 1.460 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.420 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 7.040 0.785 8.845 1.005 ;
        RECT 11.495 0.785 12.415 1.015 ;
        RECT 0.005 0.105 12.415 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.610 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 12.420 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 11.995 1.495 12.335 2.450 ;
        RECT 12.145 0.825 12.335 1.495 ;
        RECT 11.995 0.275 12.335 0.825 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 12.420 2.805 ;
        RECT 0.085 2.025 0.345 2.465 ;
        RECT 0.515 2.195 0.785 2.635 ;
        RECT 0.955 2.255 2.045 2.465 ;
        RECT 0.955 2.025 1.125 2.255 ;
        RECT 2.270 2.085 2.520 2.465 ;
        RECT 2.690 2.140 2.985 2.635 ;
        RECT 0.085 1.845 1.125 2.025 ;
        RECT 1.295 1.845 1.695 2.085 ;
        RECT 0.540 0.765 0.820 1.675 ;
        RECT 1.505 0.710 1.695 1.845 ;
        RECT 1.865 1.770 2.520 2.085 ;
        RECT 3.255 2.000 3.425 2.325 ;
        RECT 3.595 2.275 3.925 2.635 ;
        RECT 4.095 2.135 4.440 2.465 ;
        RECT 3.255 1.990 3.985 2.000 ;
        RECT 3.255 1.830 3.995 1.990 ;
        RECT 1.865 0.905 2.200 1.770 ;
        RECT 2.370 1.075 2.700 1.600 ;
        RECT 1.865 0.715 2.520 0.905 ;
        RECT 3.735 0.885 3.995 1.830 ;
        RECT 1.505 0.705 1.675 0.710 ;
        RECT 1.495 0.665 1.675 0.705 ;
        RECT 1.475 0.660 1.675 0.665 ;
        RECT 1.475 0.645 1.670 0.660 ;
        RECT 1.460 0.635 1.665 0.645 ;
        RECT 1.445 0.630 1.665 0.635 ;
        RECT 1.440 0.620 1.665 0.630 ;
        RECT 1.430 0.615 1.660 0.620 ;
        RECT 1.420 0.610 1.660 0.615 ;
        RECT 1.405 0.605 1.660 0.610 ;
        RECT 1.395 0.600 1.660 0.605 ;
        RECT 1.380 0.595 1.660 0.600 ;
        RECT 0.085 0.085 0.700 0.595 ;
        RECT 0.870 0.575 1.650 0.595 ;
        RECT 0.870 0.555 1.640 0.575 ;
        RECT 0.870 0.255 1.625 0.555 ;
        RECT 1.825 0.085 2.090 0.545 ;
        RECT 2.260 0.255 2.520 0.715 ;
        RECT 3.270 0.715 3.995 0.885 ;
        RECT 4.165 1.420 4.440 2.135 ;
        RECT 4.615 1.615 4.830 2.465 ;
        RECT 5.035 2.135 5.755 2.465 ;
        RECT 5.945 2.275 6.330 2.635 ;
        RECT 4.615 1.590 4.915 1.615 ;
        RECT 4.660 1.445 4.915 1.590 ;
        RECT 5.205 1.575 5.415 1.955 ;
        RECT 4.165 1.090 4.490 1.420 ;
        RECT 2.690 0.085 3.100 0.555 ;
        RECT 3.270 0.255 3.455 0.715 ;
        RECT 4.165 0.585 4.335 1.090 ;
        RECT 4.660 0.920 4.830 1.445 ;
        RECT 5.585 1.395 5.755 2.135 ;
        RECT 6.605 2.105 6.820 2.450 ;
        RECT 7.060 2.125 8.015 2.635 ;
        RECT 8.185 2.125 8.990 2.460 ;
        RECT 9.160 2.235 9.490 2.635 ;
        RECT 5.925 1.935 6.820 2.105 ;
        RECT 8.820 2.065 8.990 2.125 ;
        RECT 9.660 2.065 9.965 2.450 ;
        RECT 10.155 2.235 10.485 2.635 ;
        RECT 5.925 1.575 6.095 1.935 ;
        RECT 6.640 1.445 7.065 1.765 ;
        RECT 7.235 1.670 8.135 1.955 ;
        RECT 5.085 1.275 6.475 1.395 ;
        RECT 7.355 1.275 7.715 1.325 ;
        RECT 3.625 0.085 3.955 0.545 ;
        RECT 4.125 0.255 4.335 0.585 ;
        RECT 4.505 0.255 4.830 0.920 ;
        RECT 5.000 1.225 7.715 1.275 ;
        RECT 5.000 0.255 5.440 1.225 ;
        RECT 5.645 0.805 5.975 1.015 ;
        RECT 6.305 0.975 7.715 1.225 ;
        RECT 7.885 0.905 8.135 1.670 ;
        RECT 8.425 1.075 8.650 1.905 ;
        RECT 8.820 1.895 10.485 2.065 ;
        RECT 8.880 1.545 9.945 1.725 ;
        RECT 10.155 1.605 10.485 1.895 ;
        RECT 8.880 1.425 9.135 1.545 ;
        RECT 10.655 1.365 10.915 2.465 ;
        RECT 8.820 0.905 9.105 1.255 ;
        RECT 5.645 0.635 6.535 0.805 ;
        RECT 5.610 0.085 6.095 0.465 ;
        RECT 6.285 0.255 6.535 0.635 ;
        RECT 6.705 0.085 7.715 0.805 ;
        RECT 7.885 0.720 9.105 0.905 ;
        RECT 9.320 1.195 10.915 1.365 ;
        RECT 9.320 0.855 9.530 1.195 ;
        RECT 9.710 0.785 10.515 1.015 ;
        RECT 9.710 0.545 9.910 0.785 ;
        RECT 10.685 0.585 10.915 1.195 ;
        RECT 8.465 0.275 9.910 0.545 ;
        RECT 10.115 0.085 10.365 0.545 ;
        RECT 10.575 0.255 10.915 0.585 ;
        RECT 11.085 1.325 11.345 2.465 ;
        RECT 11.515 1.790 11.825 2.635 ;
        RECT 11.085 0.995 11.975 1.325 ;
        RECT 11.085 0.255 11.345 0.995 ;
        RECT 11.515 0.085 11.825 0.825 ;
        RECT 0.000 -0.085 12.420 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 0.605 1.105 0.775 1.275 ;
        RECT 1.525 1.445 1.695 1.615 ;
        RECT 3.825 1.785 3.995 1.955 ;
        RECT 2.445 1.105 2.615 1.275 ;
        RECT 5.205 1.785 5.375 1.955 ;
        RECT 4.745 1.445 4.915 1.615 ;
        RECT 4.285 1.105 4.455 1.275 ;
        RECT 7.560 1.785 7.730 1.955 ;
        RECT 8.940 1.445 9.110 1.615 ;
        RECT 8.480 1.105 8.650 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
      LAYER met1 ;
        RECT 3.765 1.940 4.055 1.985 ;
        RECT 5.145 1.940 5.435 1.985 ;
        RECT 7.500 1.940 7.790 1.985 ;
        RECT 3.765 1.800 7.790 1.940 ;
        RECT 3.765 1.755 4.055 1.800 ;
        RECT 5.145 1.755 5.435 1.800 ;
        RECT 7.500 1.755 7.790 1.800 ;
        RECT 1.465 1.600 1.755 1.645 ;
        RECT 4.685 1.600 4.975 1.645 ;
        RECT 1.465 1.460 4.975 1.600 ;
        RECT 1.465 1.415 1.755 1.460 ;
        RECT 4.685 1.415 4.975 1.460 ;
        RECT 4.225 1.260 4.515 1.305 ;
        RECT 8.420 1.260 8.710 1.305 ;
        RECT 4.225 1.120 8.710 1.260 ;
        RECT 4.225 1.075 4.515 1.120 ;
        RECT 8.420 1.075 8.710 1.120 ;
  END
END sky130_fd_sc_hd__sdfstp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfstp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.880 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.615 3.085 1.960 ;
        RECT 2.905 1.055 3.565 1.615 ;
        RECT 2.905 0.725 3.100 1.055 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.050 0.765 1.335 1.675 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.340 1.675 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER met1 ;
        RECT 0.545 1.260 0.835 1.305 ;
        RECT 2.385 1.260 2.675 1.305 ;
        RECT 0.545 1.120 2.675 1.260 ;
        RECT 0.545 1.075 0.835 1.120 ;
        RECT 2.385 1.075 2.675 1.120 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 6.580 1.600 6.870 1.645 ;
        RECT 8.880 1.600 9.170 1.645 ;
        RECT 6.580 1.460 9.170 1.600 ;
        RECT 6.580 1.415 6.870 1.460 ;
        RECT 8.880 1.415 9.170 1.460 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 12.880 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 7.040 0.785 8.845 1.005 ;
        RECT 11.490 0.785 12.875 1.015 ;
        RECT 0.005 0.105 12.875 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 13.070 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 12.880 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.519750 ;
    PORT
      LAYER li1 ;
        RECT 12.035 1.495 12.365 2.450 ;
        RECT 12.145 0.825 12.365 1.495 ;
        RECT 12.035 0.255 12.365 0.825 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 12.880 2.805 ;
        RECT 0.085 2.025 0.345 2.465 ;
        RECT 0.515 2.195 0.785 2.635 ;
        RECT 0.955 2.255 2.045 2.465 ;
        RECT 0.955 2.025 1.125 2.255 ;
        RECT 2.270 2.085 2.520 2.465 ;
        RECT 2.690 2.140 2.985 2.635 ;
        RECT 0.085 1.845 1.125 2.025 ;
        RECT 1.295 1.845 1.695 2.085 ;
        RECT 0.540 0.765 0.820 1.675 ;
        RECT 1.505 0.710 1.695 1.845 ;
        RECT 1.865 1.770 2.520 2.085 ;
        RECT 3.255 2.000 3.425 2.325 ;
        RECT 3.595 2.275 3.925 2.635 ;
        RECT 4.095 2.135 4.440 2.465 ;
        RECT 3.255 1.990 3.985 2.000 ;
        RECT 3.255 1.830 3.995 1.990 ;
        RECT 1.865 0.905 2.200 1.770 ;
        RECT 2.370 1.075 2.700 1.600 ;
        RECT 1.865 0.715 2.520 0.905 ;
        RECT 3.735 0.885 3.995 1.830 ;
        RECT 1.505 0.705 1.675 0.710 ;
        RECT 1.495 0.665 1.675 0.705 ;
        RECT 1.475 0.660 1.675 0.665 ;
        RECT 1.475 0.645 1.670 0.660 ;
        RECT 1.460 0.635 1.665 0.645 ;
        RECT 1.445 0.630 1.665 0.635 ;
        RECT 1.440 0.620 1.665 0.630 ;
        RECT 1.430 0.615 1.660 0.620 ;
        RECT 1.420 0.610 1.660 0.615 ;
        RECT 1.405 0.605 1.660 0.610 ;
        RECT 1.395 0.600 1.660 0.605 ;
        RECT 1.380 0.595 1.660 0.600 ;
        RECT 0.085 0.085 0.700 0.595 ;
        RECT 0.870 0.575 1.650 0.595 ;
        RECT 0.870 0.555 1.640 0.575 ;
        RECT 0.870 0.255 1.625 0.555 ;
        RECT 1.825 0.085 2.090 0.545 ;
        RECT 2.260 0.255 2.520 0.715 ;
        RECT 3.270 0.715 3.995 0.885 ;
        RECT 4.165 1.420 4.440 2.135 ;
        RECT 4.615 1.615 4.830 2.465 ;
        RECT 5.035 2.135 5.755 2.465 ;
        RECT 5.945 2.275 6.330 2.635 ;
        RECT 4.615 1.590 4.915 1.615 ;
        RECT 4.660 1.445 4.915 1.590 ;
        RECT 5.205 1.575 5.415 1.955 ;
        RECT 4.165 1.090 4.490 1.420 ;
        RECT 2.690 0.085 3.100 0.555 ;
        RECT 3.270 0.255 3.455 0.715 ;
        RECT 4.165 0.585 4.335 1.090 ;
        RECT 4.660 0.920 4.830 1.445 ;
        RECT 5.585 1.395 5.755 2.135 ;
        RECT 6.605 2.105 6.820 2.450 ;
        RECT 7.060 2.125 8.015 2.635 ;
        RECT 8.185 2.125 8.990 2.460 ;
        RECT 9.160 2.235 9.490 2.635 ;
        RECT 5.925 1.935 6.820 2.105 ;
        RECT 8.820 2.065 8.990 2.125 ;
        RECT 9.660 2.065 9.965 2.450 ;
        RECT 10.155 2.235 10.485 2.635 ;
        RECT 5.925 1.575 6.095 1.935 ;
        RECT 6.640 1.445 7.065 1.765 ;
        RECT 7.235 1.670 8.135 1.955 ;
        RECT 5.085 1.275 6.475 1.395 ;
        RECT 7.355 1.275 7.715 1.325 ;
        RECT 3.625 0.085 3.955 0.545 ;
        RECT 4.125 0.255 4.335 0.585 ;
        RECT 4.505 0.255 4.830 0.920 ;
        RECT 5.000 1.225 7.715 1.275 ;
        RECT 5.000 0.255 5.440 1.225 ;
        RECT 5.645 0.805 5.975 1.015 ;
        RECT 6.305 0.975 7.715 1.225 ;
        RECT 7.885 0.905 8.135 1.670 ;
        RECT 8.425 1.075 8.650 1.905 ;
        RECT 8.820 1.895 10.485 2.065 ;
        RECT 8.880 1.545 9.945 1.725 ;
        RECT 10.155 1.605 10.485 1.895 ;
        RECT 8.880 1.425 9.135 1.545 ;
        RECT 10.655 1.365 10.915 2.465 ;
        RECT 8.820 0.905 9.105 1.255 ;
        RECT 5.645 0.635 6.535 0.805 ;
        RECT 5.610 0.085 6.095 0.465 ;
        RECT 6.285 0.255 6.535 0.635 ;
        RECT 6.705 0.085 7.715 0.805 ;
        RECT 7.885 0.720 9.105 0.905 ;
        RECT 9.320 1.195 10.915 1.365 ;
        RECT 9.320 0.855 9.530 1.195 ;
        RECT 9.710 0.785 10.515 1.015 ;
        RECT 9.710 0.545 9.910 0.785 ;
        RECT 10.685 0.585 10.915 1.195 ;
        RECT 8.465 0.275 9.910 0.545 ;
        RECT 10.115 0.085 10.365 0.545 ;
        RECT 10.575 0.255 10.915 0.585 ;
        RECT 11.085 1.325 11.345 2.465 ;
        RECT 11.570 1.790 11.820 2.635 ;
        RECT 12.535 1.495 12.795 2.635 ;
        RECT 11.085 0.995 11.975 1.325 ;
        RECT 11.085 0.255 11.345 0.995 ;
        RECT 11.570 0.085 11.865 0.825 ;
        RECT 12.535 0.085 12.795 0.885 ;
        RECT 0.000 -0.085 12.880 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 0.605 1.105 0.775 1.275 ;
        RECT 1.525 1.445 1.695 1.615 ;
        RECT 3.825 1.785 3.995 1.955 ;
        RECT 2.445 1.105 2.615 1.275 ;
        RECT 5.205 1.785 5.375 1.955 ;
        RECT 4.745 1.445 4.915 1.615 ;
        RECT 4.285 1.105 4.455 1.275 ;
        RECT 7.560 1.785 7.730 1.955 ;
        RECT 8.940 1.445 9.110 1.615 ;
        RECT 8.480 1.105 8.650 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
      LAYER met1 ;
        RECT 3.765 1.940 4.055 1.985 ;
        RECT 5.145 1.940 5.435 1.985 ;
        RECT 7.500 1.940 7.790 1.985 ;
        RECT 3.765 1.800 7.790 1.940 ;
        RECT 3.765 1.755 4.055 1.800 ;
        RECT 5.145 1.755 5.435 1.800 ;
        RECT 7.500 1.755 7.790 1.800 ;
        RECT 1.465 1.600 1.755 1.645 ;
        RECT 4.685 1.600 4.975 1.645 ;
        RECT 1.465 1.460 4.975 1.600 ;
        RECT 1.465 1.415 1.755 1.460 ;
        RECT 4.685 1.415 4.975 1.460 ;
        RECT 4.225 1.260 4.515 1.305 ;
        RECT 8.420 1.260 8.710 1.305 ;
        RECT 4.225 1.120 8.710 1.260 ;
        RECT 4.225 1.075 4.515 1.120 ;
        RECT 8.420 1.075 8.710 1.120 ;
  END
END sky130_fd_sc_hd__sdfstp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfstp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfstp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.800 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.905 1.615 3.085 1.960 ;
        RECT 2.905 1.055 3.565 1.615 ;
        RECT 2.905 0.725 3.100 1.055 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.050 0.765 1.335 1.675 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.765 0.340 1.675 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER met1 ;
        RECT 0.545 1.260 0.835 1.305 ;
        RECT 2.385 1.260 2.675 1.305 ;
        RECT 0.545 1.120 2.675 1.260 ;
        RECT 0.545 1.075 0.835 1.120 ;
        RECT 2.385 1.075 2.675 1.120 ;
    END
  END SCE
  PIN SET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met1 ;
        RECT 6.580 1.600 6.870 1.645 ;
        RECT 8.880 1.600 9.170 1.645 ;
        RECT 6.580 1.460 9.170 1.600 ;
        RECT 6.580 1.415 6.870 1.460 ;
        RECT 8.880 1.415 9.170 1.460 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 13.800 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 7.040 0.785 8.845 1.005 ;
        RECT 11.005 0.785 13.720 1.015 ;
        RECT 0.005 0.105 13.720 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 13.990 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 13.800 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 12.040 1.495 12.370 2.450 ;
        RECT 12.145 1.325 12.370 1.495 ;
        RECT 12.880 1.325 13.210 2.465 ;
        RECT 12.145 1.055 13.210 1.325 ;
        RECT 12.145 0.825 12.370 1.055 ;
        RECT 12.040 0.275 12.370 0.825 ;
        RECT 12.880 0.255 13.210 1.055 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 13.800 2.805 ;
        RECT 0.085 2.025 0.345 2.465 ;
        RECT 0.515 2.195 0.785 2.635 ;
        RECT 0.955 2.255 2.045 2.465 ;
        RECT 0.955 2.025 1.125 2.255 ;
        RECT 2.270 2.085 2.520 2.465 ;
        RECT 2.690 2.140 2.985 2.635 ;
        RECT 0.085 1.845 1.125 2.025 ;
        RECT 1.295 1.845 1.695 2.085 ;
        RECT 0.540 0.765 0.820 1.675 ;
        RECT 1.505 0.710 1.695 1.845 ;
        RECT 1.865 1.770 2.520 2.085 ;
        RECT 3.255 2.000 3.425 2.325 ;
        RECT 3.595 2.275 3.925 2.635 ;
        RECT 4.095 2.135 4.440 2.465 ;
        RECT 3.255 1.990 3.985 2.000 ;
        RECT 3.255 1.830 3.995 1.990 ;
        RECT 1.865 0.905 2.200 1.770 ;
        RECT 2.370 1.075 2.700 1.600 ;
        RECT 1.865 0.715 2.520 0.905 ;
        RECT 3.735 0.885 3.995 1.830 ;
        RECT 1.505 0.705 1.675 0.710 ;
        RECT 1.495 0.665 1.675 0.705 ;
        RECT 1.475 0.660 1.675 0.665 ;
        RECT 1.475 0.645 1.670 0.660 ;
        RECT 1.460 0.635 1.665 0.645 ;
        RECT 1.445 0.630 1.665 0.635 ;
        RECT 1.440 0.620 1.665 0.630 ;
        RECT 1.430 0.615 1.660 0.620 ;
        RECT 1.420 0.610 1.660 0.615 ;
        RECT 1.405 0.605 1.660 0.610 ;
        RECT 1.395 0.600 1.660 0.605 ;
        RECT 1.380 0.595 1.660 0.600 ;
        RECT 0.085 0.085 0.700 0.595 ;
        RECT 0.870 0.575 1.650 0.595 ;
        RECT 0.870 0.555 1.640 0.575 ;
        RECT 0.870 0.255 1.625 0.555 ;
        RECT 1.825 0.085 2.090 0.545 ;
        RECT 2.260 0.255 2.520 0.715 ;
        RECT 3.270 0.715 3.995 0.885 ;
        RECT 4.165 1.420 4.440 2.135 ;
        RECT 4.615 1.615 4.830 2.465 ;
        RECT 5.035 2.135 5.755 2.465 ;
        RECT 5.945 2.275 6.330 2.635 ;
        RECT 4.615 1.590 4.915 1.615 ;
        RECT 4.660 1.445 4.915 1.590 ;
        RECT 5.205 1.575 5.415 1.955 ;
        RECT 4.165 1.090 4.490 1.420 ;
        RECT 2.690 0.085 3.100 0.555 ;
        RECT 3.270 0.255 3.455 0.715 ;
        RECT 4.165 0.585 4.335 1.090 ;
        RECT 4.660 0.920 4.830 1.445 ;
        RECT 5.585 1.395 5.755 2.135 ;
        RECT 6.605 2.105 6.820 2.450 ;
        RECT 7.060 2.125 8.015 2.635 ;
        RECT 8.185 2.125 8.990 2.460 ;
        RECT 9.160 2.235 9.490 2.635 ;
        RECT 5.925 1.935 6.820 2.105 ;
        RECT 8.820 2.065 8.990 2.125 ;
        RECT 9.660 2.065 9.965 2.450 ;
        RECT 10.155 2.235 10.485 2.635 ;
        RECT 5.925 1.575 6.095 1.935 ;
        RECT 6.640 1.445 7.065 1.765 ;
        RECT 7.235 1.670 8.135 1.955 ;
        RECT 5.085 1.275 6.475 1.395 ;
        RECT 7.355 1.275 7.715 1.325 ;
        RECT 3.625 0.085 3.955 0.545 ;
        RECT 4.125 0.255 4.335 0.585 ;
        RECT 4.505 0.255 4.830 0.920 ;
        RECT 5.000 1.225 7.715 1.275 ;
        RECT 5.000 0.255 5.440 1.225 ;
        RECT 5.645 0.805 5.975 1.015 ;
        RECT 6.305 0.975 7.715 1.225 ;
        RECT 7.885 0.905 8.135 1.670 ;
        RECT 8.425 1.075 8.650 1.905 ;
        RECT 8.820 1.895 10.485 2.065 ;
        RECT 8.880 1.545 9.945 1.725 ;
        RECT 10.155 1.605 10.485 1.895 ;
        RECT 8.880 1.425 9.135 1.545 ;
        RECT 10.655 1.365 10.915 2.465 ;
        RECT 8.820 0.905 9.105 1.255 ;
        RECT 5.645 0.635 6.535 0.805 ;
        RECT 5.610 0.085 6.095 0.465 ;
        RECT 6.285 0.255 6.535 0.635 ;
        RECT 6.705 0.085 7.715 0.805 ;
        RECT 7.885 0.720 9.105 0.905 ;
        RECT 9.320 1.195 10.915 1.365 ;
        RECT 9.320 0.855 9.530 1.195 ;
        RECT 9.710 0.785 10.515 1.015 ;
        RECT 9.710 0.545 9.910 0.785 ;
        RECT 10.685 0.585 10.915 1.195 ;
        RECT 8.465 0.275 9.910 0.545 ;
        RECT 10.115 0.085 10.365 0.545 ;
        RECT 10.575 0.255 10.915 0.585 ;
        RECT 11.085 1.325 11.345 2.465 ;
        RECT 11.515 1.495 11.870 2.635 ;
        RECT 12.540 1.495 12.710 2.635 ;
        RECT 13.380 1.495 13.715 2.635 ;
        RECT 11.085 0.995 11.975 1.325 ;
        RECT 11.085 0.255 11.345 0.995 ;
        RECT 11.515 0.085 11.870 0.825 ;
        RECT 12.540 0.085 12.710 0.885 ;
        RECT 13.380 0.085 13.715 0.885 ;
        RECT 0.000 -0.085 13.800 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 0.605 1.105 0.775 1.275 ;
        RECT 1.525 1.445 1.695 1.615 ;
        RECT 3.825 1.785 3.995 1.955 ;
        RECT 2.445 1.105 2.615 1.275 ;
        RECT 5.205 1.785 5.375 1.955 ;
        RECT 4.745 1.445 4.915 1.615 ;
        RECT 4.285 1.105 4.455 1.275 ;
        RECT 7.560 1.785 7.730 1.955 ;
        RECT 8.940 1.445 9.110 1.615 ;
        RECT 8.480 1.105 8.650 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
      LAYER met1 ;
        RECT 3.765 1.940 4.055 1.985 ;
        RECT 5.145 1.940 5.435 1.985 ;
        RECT 7.500 1.940 7.790 1.985 ;
        RECT 3.765 1.800 7.790 1.940 ;
        RECT 3.765 1.755 4.055 1.800 ;
        RECT 5.145 1.755 5.435 1.800 ;
        RECT 7.500 1.755 7.790 1.800 ;
        RECT 1.465 1.600 1.755 1.645 ;
        RECT 4.685 1.600 4.975 1.645 ;
        RECT 1.465 1.460 4.975 1.600 ;
        RECT 1.465 1.415 1.755 1.460 ;
        RECT 4.685 1.415 4.975 1.460 ;
        RECT 4.225 1.260 4.515 1.305 ;
        RECT 8.420 1.260 8.710 1.305 ;
        RECT 4.225 1.120 8.710 1.260 ;
        RECT 4.225 1.075 4.515 1.120 ;
        RECT 8.420 1.075 8.710 1.120 ;
  END
END sky130_fd_sc_hd__sdfstp_4

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.440 1.355 2.775 1.685 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 3.515 1.055 3.995 1.655 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 1.760 0.880 1.930 1.685 ;
        RECT 1.760 0.875 1.940 0.880 ;
        RECT 1.760 0.870 1.945 0.875 ;
        RECT 1.760 0.860 1.950 0.870 ;
        RECT 1.760 0.855 1.955 0.860 ;
        RECT 1.760 0.850 1.960 0.855 ;
        RECT 1.760 0.840 1.965 0.850 ;
        RECT 1.760 0.835 1.970 0.840 ;
        RECT 1.760 0.820 1.975 0.835 ;
        RECT 1.760 0.810 1.990 0.820 ;
        RECT 1.760 0.785 2.010 0.810 ;
        RECT 3.065 0.785 3.235 1.115 ;
        RECT 1.760 0.750 3.235 0.785 ;
        RECT 1.790 0.735 3.235 0.750 ;
        RECT 1.805 0.725 3.235 0.735 ;
        RECT 1.820 0.715 3.235 0.725 ;
        RECT 1.830 0.705 3.235 0.715 ;
        RECT 1.840 0.690 3.235 0.705 ;
        RECT 1.860 0.655 3.235 0.690 ;
        RECT 1.875 0.615 3.235 0.655 ;
        RECT 2.455 0.305 2.630 0.615 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.825 0.785 6.735 1.005 ;
        RECT 8.250 0.785 11.025 1.015 ;
        RECT 0.005 0.725 4.085 0.785 ;
        RECT 5.095 0.725 11.025 0.785 ;
        RECT 0.005 0.105 11.025 0.725 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 9.200 1.540 9.530 2.465 ;
        RECT 9.200 1.505 9.610 1.540 ;
        RECT 9.355 1.430 9.610 1.505 ;
        RECT 9.390 0.825 9.610 1.430 ;
        RECT 9.180 0.790 9.610 0.825 ;
        RECT 9.180 0.725 9.560 0.790 ;
        RECT 9.180 0.305 9.530 0.725 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 10.685 1.445 10.940 2.325 ;
        RECT 10.730 0.795 10.940 1.445 ;
        RECT 10.685 0.265 10.940 0.795 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.845 1.965 ;
        RECT 0.615 0.970 0.845 1.795 ;
        RECT 0.615 0.805 0.810 0.970 ;
        RECT 0.175 0.635 0.810 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 2.465 ;
        RECT 1.420 2.075 1.705 2.445 ;
        RECT 1.875 2.245 2.205 2.635 ;
        RECT 2.675 2.245 3.570 2.415 ;
        RECT 1.420 1.860 3.230 2.075 ;
        RECT 1.420 0.585 1.590 1.860 ;
        RECT 2.100 1.125 2.270 1.860 ;
        RECT 3.060 1.685 3.230 1.860 ;
        RECT 3.400 1.995 3.570 2.245 ;
        RECT 3.740 2.165 3.910 2.635 ;
        RECT 4.165 2.070 4.450 2.440 ;
        RECT 4.645 2.190 5.715 2.360 ;
        RECT 4.165 1.995 4.335 2.070 ;
        RECT 3.400 1.825 4.335 1.995 ;
        RECT 3.060 1.355 3.255 1.685 ;
        RECT 2.100 0.955 2.445 1.125 ;
        RECT 4.165 0.885 4.335 1.825 ;
        RECT 3.405 0.715 4.335 0.885 ;
        RECT 1.420 0.255 1.705 0.585 ;
        RECT 3.405 0.445 3.575 0.715 ;
        RECT 1.955 0.085 2.285 0.445 ;
        RECT 2.800 0.275 3.575 0.445 ;
        RECT 3.745 0.085 3.945 0.545 ;
        RECT 4.165 0.535 4.335 0.715 ;
        RECT 4.505 1.035 4.745 1.905 ;
        RECT 4.935 1.655 5.375 2.010 ;
        RECT 5.545 1.575 5.715 2.190 ;
        RECT 5.885 1.835 6.055 2.635 ;
        RECT 6.225 2.135 6.475 2.465 ;
        RECT 6.700 2.165 7.585 2.335 ;
        RECT 5.545 1.485 6.055 1.575 ;
        RECT 5.255 1.315 6.055 1.485 ;
        RECT 4.505 0.705 5.085 1.035 ;
        RECT 5.255 0.535 5.425 1.315 ;
        RECT 5.885 1.245 6.055 1.315 ;
        RECT 5.595 1.065 5.765 1.095 ;
        RECT 6.225 1.065 6.395 2.135 ;
        RECT 6.565 1.245 6.755 1.965 ;
        RECT 6.925 1.575 7.245 1.905 ;
        RECT 5.595 0.765 6.395 1.065 ;
        RECT 6.925 1.035 7.115 1.575 ;
        RECT 7.415 1.405 7.585 2.165 ;
        RECT 7.765 2.135 8.070 2.635 ;
        RECT 8.380 1.905 8.670 2.455 ;
        RECT 7.755 1.575 8.670 1.905 ;
        RECT 8.840 1.625 9.010 2.635 ;
        RECT 9.700 1.685 10.030 2.425 ;
        RECT 4.165 0.365 4.515 0.535 ;
        RECT 4.685 0.365 5.425 0.535 ;
        RECT 5.675 0.085 6.045 0.585 ;
        RECT 6.225 0.535 6.395 0.765 ;
        RECT 6.565 0.705 7.115 1.035 ;
        RECT 7.285 1.325 7.585 1.405 ;
        RECT 8.485 1.325 8.670 1.575 ;
        RECT 9.780 1.325 10.030 1.685 ;
        RECT 10.210 1.495 10.515 2.635 ;
        RECT 7.285 0.995 8.315 1.325 ;
        RECT 8.485 0.995 9.220 1.325 ;
        RECT 9.780 0.995 10.560 1.325 ;
        RECT 7.285 0.535 7.455 0.995 ;
        RECT 8.485 0.825 8.670 0.995 ;
        RECT 6.225 0.365 6.685 0.535 ;
        RECT 6.915 0.365 7.455 0.535 ;
        RECT 7.700 0.085 8.070 0.615 ;
        RECT 8.340 0.300 8.670 0.825 ;
        RECT 8.840 0.085 9.010 0.695 ;
        RECT 9.780 0.620 9.950 0.995 ;
        RECT 9.700 0.345 9.950 0.620 ;
        RECT 10.185 0.085 10.515 0.805 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 0.645 1.785 0.815 1.955 ;
        RECT 1.015 0.765 1.185 0.935 ;
        RECT 5.165 1.785 5.335 1.955 ;
        RECT 4.745 0.765 4.915 0.935 ;
        RECT 6.575 1.785 6.745 1.955 ;
        RECT 6.585 0.765 6.755 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
      LAYER met1 ;
        RECT 0.585 1.940 0.875 1.985 ;
        RECT 5.105 1.940 5.395 1.985 ;
        RECT 6.515 1.940 6.805 1.985 ;
        RECT 0.585 1.800 6.805 1.940 ;
        RECT 0.585 1.755 0.875 1.800 ;
        RECT 5.105 1.755 5.395 1.800 ;
        RECT 6.515 1.755 6.805 1.800 ;
        RECT 0.955 0.920 1.245 0.965 ;
        RECT 4.685 0.920 4.975 0.965 ;
        RECT 6.525 0.920 6.815 0.965 ;
        RECT 0.955 0.780 6.815 0.920 ;
        RECT 0.955 0.735 1.245 0.780 ;
        RECT 4.685 0.735 4.975 0.780 ;
        RECT 6.525 0.735 6.815 0.780 ;
  END
END sky130_fd_sc_hd__sdfxbp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.960 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.460 1.355 2.795 1.685 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 3.535 1.035 4.035 1.655 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 1.780 0.785 1.950 1.685 ;
        RECT 3.085 0.785 3.255 1.115 ;
        RECT 1.780 0.615 3.255 0.785 ;
        RECT 2.475 0.305 2.650 0.615 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.960 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.865 0.785 6.775 1.005 ;
        RECT 8.305 0.785 11.950 1.015 ;
        RECT 0.005 0.725 4.125 0.785 ;
        RECT 5.135 0.725 11.950 0.785 ;
        RECT 0.005 0.105 11.950 0.725 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 12.150 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.960 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 9.255 1.530 9.585 2.430 ;
        RECT 9.255 1.495 9.615 1.530 ;
        RECT 9.410 1.430 9.615 1.495 ;
        RECT 9.445 0.890 9.615 1.430 ;
        RECT 9.410 0.825 9.615 0.890 ;
        RECT 9.255 0.790 9.615 0.825 ;
        RECT 9.255 0.255 9.585 0.790 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 11.190 1.445 11.440 2.325 ;
        RECT 11.235 0.795 11.440 1.445 ;
        RECT 11.190 0.265 11.440 0.795 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.960 2.805 ;
        RECT 0.180 1.965 0.350 2.465 ;
        RECT 0.520 2.135 0.850 2.635 ;
        RECT 0.180 1.795 0.845 1.965 ;
        RECT 0.615 0.970 0.845 1.795 ;
        RECT 0.615 0.805 0.810 0.970 ;
        RECT 0.175 0.635 0.810 0.805 ;
        RECT 1.020 0.715 1.245 2.465 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.245 0.715 ;
        RECT 1.435 2.075 1.710 2.445 ;
        RECT 1.880 2.245 2.210 2.635 ;
        RECT 2.695 2.245 3.590 2.415 ;
        RECT 1.435 1.860 3.250 2.075 ;
        RECT 1.435 0.445 1.605 1.860 ;
        RECT 2.120 1.125 2.290 1.860 ;
        RECT 3.080 1.685 3.250 1.860 ;
        RECT 3.420 1.995 3.590 2.245 ;
        RECT 3.760 2.165 3.930 2.635 ;
        RECT 4.205 2.065 4.485 2.440 ;
        RECT 4.685 2.190 5.755 2.360 ;
        RECT 4.205 1.995 4.375 2.065 ;
        RECT 3.420 1.825 4.375 1.995 ;
        RECT 3.080 1.355 3.275 1.685 ;
        RECT 2.120 0.955 2.465 1.125 ;
        RECT 4.205 0.865 4.375 1.825 ;
        RECT 3.425 0.695 4.375 0.865 ;
        RECT 4.545 1.035 4.785 1.905 ;
        RECT 4.975 1.655 5.415 2.010 ;
        RECT 5.585 1.575 5.755 2.190 ;
        RECT 5.925 1.835 6.095 2.635 ;
        RECT 6.265 2.135 6.515 2.465 ;
        RECT 6.740 2.165 7.625 2.335 ;
        RECT 5.585 1.485 6.095 1.575 ;
        RECT 5.295 1.315 6.095 1.485 ;
        RECT 4.545 0.705 5.125 1.035 ;
        RECT 3.425 0.445 3.595 0.695 ;
        RECT 4.205 0.535 4.375 0.695 ;
        RECT 5.295 0.535 5.465 1.315 ;
        RECT 5.925 1.245 6.095 1.315 ;
        RECT 5.635 1.065 5.805 1.095 ;
        RECT 6.265 1.065 6.435 2.135 ;
        RECT 6.605 1.245 6.795 1.965 ;
        RECT 6.965 1.575 7.285 1.905 ;
        RECT 5.635 0.765 6.435 1.065 ;
        RECT 6.965 1.035 7.155 1.575 ;
        RECT 7.455 1.405 7.625 2.165 ;
        RECT 7.805 2.135 8.110 2.635 ;
        RECT 8.395 1.905 8.725 2.455 ;
        RECT 7.795 1.575 8.725 1.905 ;
        RECT 8.895 1.625 9.075 2.635 ;
        RECT 9.765 1.615 9.935 2.635 ;
        RECT 1.435 0.275 1.805 0.445 ;
        RECT 1.975 0.085 2.305 0.445 ;
        RECT 2.820 0.275 3.595 0.445 ;
        RECT 3.765 0.085 3.965 0.525 ;
        RECT 4.205 0.365 4.555 0.535 ;
        RECT 4.725 0.365 5.465 0.535 ;
        RECT 5.715 0.085 6.085 0.585 ;
        RECT 6.265 0.535 6.435 0.765 ;
        RECT 6.605 0.705 7.155 1.035 ;
        RECT 7.325 1.325 7.625 1.405 ;
        RECT 8.540 1.325 8.725 1.575 ;
        RECT 10.205 1.325 10.535 2.425 ;
        RECT 10.715 1.495 11.020 2.635 ;
        RECT 11.610 1.395 11.780 2.635 ;
        RECT 7.325 0.995 8.370 1.325 ;
        RECT 8.540 0.995 9.275 1.325 ;
        RECT 10.205 0.995 11.065 1.325 ;
        RECT 7.325 0.535 7.495 0.995 ;
        RECT 8.540 0.825 8.725 0.995 ;
        RECT 6.265 0.365 6.725 0.535 ;
        RECT 6.955 0.365 7.495 0.535 ;
        RECT 7.740 0.085 8.110 0.615 ;
        RECT 8.360 0.300 8.725 0.825 ;
        RECT 8.895 0.085 9.085 0.695 ;
        RECT 9.755 0.085 9.985 0.690 ;
        RECT 10.205 0.345 10.455 0.995 ;
        RECT 10.690 0.085 11.020 0.805 ;
        RECT 11.610 0.085 11.780 0.955 ;
        RECT 0.000 -0.085 11.960 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 0.645 1.785 0.815 1.955 ;
        RECT 1.050 0.765 1.220 0.935 ;
        RECT 5.205 1.785 5.375 1.955 ;
        RECT 4.745 0.765 4.915 0.935 ;
        RECT 6.625 1.785 6.795 1.955 ;
        RECT 6.640 0.765 6.810 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
      LAYER met1 ;
        RECT 0.585 1.940 0.875 1.985 ;
        RECT 5.145 1.940 5.435 1.985 ;
        RECT 6.565 1.940 6.855 1.985 ;
        RECT 0.585 1.800 6.855 1.940 ;
        RECT 0.585 1.755 0.875 1.800 ;
        RECT 5.145 1.755 5.435 1.800 ;
        RECT 6.565 1.755 6.855 1.800 ;
        RECT 0.990 0.920 1.280 0.965 ;
        RECT 4.685 0.920 4.975 0.965 ;
        RECT 6.580 0.920 6.870 0.965 ;
        RECT 0.990 0.780 6.870 0.920 ;
        RECT 0.990 0.735 1.280 0.780 ;
        RECT 4.685 0.735 4.975 0.780 ;
        RECT 6.580 0.735 6.870 0.780 ;
  END
END sky130_fd_sc_hd__sdfxbp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.460 1.355 2.790 1.685 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 3.530 1.055 3.990 1.655 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 1.760 0.835 1.930 1.685 ;
        RECT 1.760 0.785 1.990 0.835 ;
        RECT 3.065 0.785 3.250 1.095 ;
        RECT 1.760 0.635 3.250 0.785 ;
        RECT 1.870 0.615 3.250 0.635 ;
        RECT 2.475 0.305 2.650 0.615 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.840 0.785 6.750 1.005 ;
        RECT 8.265 0.785 9.650 1.015 ;
        RECT 0.005 0.725 4.105 0.785 ;
        RECT 5.110 0.725 9.650 0.785 ;
        RECT 0.005 0.105 9.650 0.725 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 9.230 1.505 9.575 2.395 ;
        RECT 9.405 0.820 9.575 1.505 ;
        RECT 9.230 0.305 9.575 0.820 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.180 1.965 0.350 2.465 ;
        RECT 0.520 2.135 0.850 2.635 ;
        RECT 0.180 1.795 0.845 1.965 ;
        RECT 0.615 0.970 0.845 1.795 ;
        RECT 0.615 0.805 0.810 0.970 ;
        RECT 0.175 0.635 0.810 0.805 ;
        RECT 1.020 0.715 1.230 2.465 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.230 0.715 ;
        RECT 1.420 2.075 1.710 2.445 ;
        RECT 1.880 2.245 2.210 2.635 ;
        RECT 2.690 2.245 3.560 2.415 ;
        RECT 1.420 1.860 3.220 2.075 ;
        RECT 1.420 0.465 1.590 1.860 ;
        RECT 2.115 1.130 2.290 1.860 ;
        RECT 3.050 1.635 3.220 1.860 ;
        RECT 3.390 1.995 3.560 2.245 ;
        RECT 3.730 2.165 3.925 2.635 ;
        RECT 4.180 2.065 4.420 2.440 ;
        RECT 4.660 2.190 5.730 2.360 ;
        RECT 4.180 1.995 4.350 2.065 ;
        RECT 3.390 1.825 4.350 1.995 ;
        RECT 3.050 1.305 3.270 1.635 ;
        RECT 2.115 0.960 2.460 1.130 ;
        RECT 4.180 0.885 4.350 1.825 ;
        RECT 3.420 0.715 4.350 0.885 ;
        RECT 4.520 1.035 4.760 1.905 ;
        RECT 4.950 1.655 5.390 2.010 ;
        RECT 5.560 1.575 5.730 2.190 ;
        RECT 5.900 1.835 6.070 2.635 ;
        RECT 6.240 2.135 6.490 2.465 ;
        RECT 6.715 2.165 7.600 2.335 ;
        RECT 5.560 1.485 6.070 1.575 ;
        RECT 5.270 1.315 6.070 1.485 ;
        RECT 4.520 0.780 5.100 1.035 ;
        RECT 1.420 0.260 1.790 0.465 ;
        RECT 3.420 0.445 3.590 0.715 ;
        RECT 4.180 0.615 4.350 0.715 ;
        RECT 4.630 0.705 5.100 0.780 ;
        RECT 1.960 0.085 2.305 0.445 ;
        RECT 2.820 0.275 3.590 0.445 ;
        RECT 3.760 0.085 3.960 0.545 ;
        RECT 4.180 0.285 4.460 0.615 ;
        RECT 5.270 0.535 5.440 1.315 ;
        RECT 5.900 1.245 6.070 1.315 ;
        RECT 5.610 1.065 5.780 1.095 ;
        RECT 6.240 1.065 6.410 2.135 ;
        RECT 6.580 1.245 6.770 1.965 ;
        RECT 6.940 1.575 7.260 1.905 ;
        RECT 5.610 0.765 6.410 1.065 ;
        RECT 6.940 1.035 7.130 1.575 ;
        RECT 7.430 1.405 7.600 2.165 ;
        RECT 7.790 2.135 8.095 2.635 ;
        RECT 8.435 1.905 8.705 2.455 ;
        RECT 7.770 1.575 8.705 1.905 ;
        RECT 8.875 1.625 9.045 2.635 ;
        RECT 4.700 0.365 5.440 0.535 ;
        RECT 5.690 0.085 6.060 0.585 ;
        RECT 6.240 0.535 6.410 0.765 ;
        RECT 6.580 0.705 7.130 1.035 ;
        RECT 7.300 1.325 7.600 1.405 ;
        RECT 8.535 1.325 8.705 1.575 ;
        RECT 7.300 0.995 8.365 1.325 ;
        RECT 8.535 0.995 9.235 1.325 ;
        RECT 7.300 0.535 7.470 0.995 ;
        RECT 8.535 0.825 8.705 0.995 ;
        RECT 6.240 0.365 6.700 0.535 ;
        RECT 6.930 0.365 7.470 0.535 ;
        RECT 7.715 0.085 8.085 0.615 ;
        RECT 8.355 0.300 8.705 0.825 ;
        RECT 8.875 0.085 9.045 0.695 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 0.640 1.785 0.810 1.955 ;
        RECT 1.040 0.765 1.210 0.935 ;
        RECT 5.205 1.785 5.375 1.955 ;
        RECT 4.745 0.765 4.915 0.935 ;
        RECT 6.590 1.785 6.760 1.955 ;
        RECT 6.630 0.765 6.800 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 0.580 1.940 0.870 1.985 ;
        RECT 5.145 1.940 5.435 1.985 ;
        RECT 6.530 1.940 6.820 1.985 ;
        RECT 0.580 1.800 6.820 1.940 ;
        RECT 0.580 1.755 0.870 1.800 ;
        RECT 5.145 1.755 5.435 1.800 ;
        RECT 6.530 1.755 6.820 1.800 ;
        RECT 0.980 0.920 1.270 0.965 ;
        RECT 4.685 0.920 4.975 0.965 ;
        RECT 6.570 0.920 6.860 0.965 ;
        RECT 0.980 0.780 6.860 0.920 ;
        RECT 0.980 0.735 1.270 0.780 ;
        RECT 4.685 0.735 4.975 0.780 ;
        RECT 6.570 0.735 6.860 0.780 ;
  END
END sky130_fd_sc_hd__sdfxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.460 1.355 2.790 1.685 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 3.530 1.035 4.020 1.655 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 1.780 0.785 1.950 1.685 ;
        RECT 3.080 0.785 3.250 1.115 ;
        RECT 1.780 0.615 3.250 0.785 ;
        RECT 2.475 0.305 2.650 0.615 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.870 0.785 6.780 1.005 ;
        RECT 8.295 0.785 10.115 1.015 ;
        RECT 0.005 0.725 4.120 0.785 ;
        RECT 5.140 0.725 10.115 0.785 ;
        RECT 0.005 0.105 10.115 0.725 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 9.260 1.505 9.605 2.395 ;
        RECT 9.435 0.820 9.605 1.505 ;
        RECT 9.260 0.305 9.605 0.820 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.180 1.965 0.350 2.465 ;
        RECT 0.520 2.135 0.850 2.635 ;
        RECT 0.180 1.795 0.845 1.965 ;
        RECT 0.615 0.970 0.845 1.795 ;
        RECT 0.615 0.805 0.810 0.970 ;
        RECT 0.175 0.635 0.810 0.805 ;
        RECT 1.020 0.715 1.245 2.465 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.245 0.715 ;
        RECT 1.435 2.075 1.710 2.445 ;
        RECT 1.880 2.245 2.210 2.635 ;
        RECT 2.690 2.245 3.585 2.415 ;
        RECT 1.435 1.860 3.245 2.075 ;
        RECT 1.435 0.445 1.605 1.860 ;
        RECT 2.120 1.125 2.290 1.860 ;
        RECT 3.075 1.685 3.245 1.860 ;
        RECT 3.415 1.995 3.585 2.245 ;
        RECT 3.755 2.165 3.925 2.635 ;
        RECT 4.210 2.065 4.445 2.440 ;
        RECT 4.690 2.190 5.760 2.360 ;
        RECT 4.210 1.995 4.380 2.065 ;
        RECT 3.415 1.825 4.380 1.995 ;
        RECT 3.075 1.355 3.270 1.685 ;
        RECT 2.120 0.955 2.460 1.125 ;
        RECT 4.210 0.865 4.380 1.825 ;
        RECT 3.420 0.695 4.380 0.865 ;
        RECT 4.550 1.035 4.790 1.905 ;
        RECT 4.980 1.655 5.420 2.010 ;
        RECT 5.590 1.575 5.760 2.190 ;
        RECT 5.930 1.835 6.100 2.635 ;
        RECT 6.270 2.135 6.520 2.465 ;
        RECT 6.745 2.165 7.630 2.335 ;
        RECT 5.590 1.485 6.100 1.575 ;
        RECT 5.300 1.315 6.100 1.485 ;
        RECT 4.550 0.705 5.130 1.035 ;
        RECT 3.420 0.445 3.590 0.695 ;
        RECT 4.210 0.535 4.380 0.695 ;
        RECT 5.300 0.535 5.470 1.315 ;
        RECT 5.930 1.245 6.100 1.315 ;
        RECT 5.640 1.065 5.810 1.095 ;
        RECT 6.270 1.065 6.440 2.135 ;
        RECT 6.610 1.245 6.800 1.965 ;
        RECT 6.970 1.575 7.290 1.905 ;
        RECT 5.640 0.765 6.440 1.065 ;
        RECT 6.970 1.035 7.160 1.575 ;
        RECT 7.460 1.405 7.630 2.165 ;
        RECT 7.810 2.135 8.115 2.635 ;
        RECT 8.465 1.905 8.735 2.455 ;
        RECT 7.800 1.575 8.735 1.905 ;
        RECT 8.905 1.625 9.080 2.635 ;
        RECT 1.435 0.275 1.805 0.445 ;
        RECT 1.975 0.085 2.305 0.445 ;
        RECT 2.820 0.275 3.590 0.445 ;
        RECT 3.760 0.085 3.960 0.525 ;
        RECT 4.210 0.365 4.560 0.535 ;
        RECT 4.730 0.365 5.470 0.535 ;
        RECT 5.720 0.085 6.090 0.585 ;
        RECT 6.270 0.535 6.440 0.765 ;
        RECT 6.610 0.705 7.160 1.035 ;
        RECT 7.330 1.325 7.630 1.405 ;
        RECT 8.565 1.325 8.735 1.575 ;
        RECT 9.775 1.405 9.945 2.635 ;
        RECT 7.330 0.995 8.395 1.325 ;
        RECT 8.565 0.995 9.265 1.325 ;
        RECT 7.330 0.535 7.500 0.995 ;
        RECT 8.565 0.825 8.735 0.995 ;
        RECT 6.270 0.365 6.730 0.535 ;
        RECT 6.960 0.365 7.500 0.535 ;
        RECT 7.745 0.085 8.115 0.615 ;
        RECT 8.385 0.300 8.735 0.825 ;
        RECT 8.905 0.085 9.075 0.695 ;
        RECT 9.775 0.085 9.945 0.930 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 0.640 1.785 0.810 1.955 ;
        RECT 1.050 0.765 1.220 0.935 ;
        RECT 5.205 1.785 5.375 1.955 ;
        RECT 4.745 0.765 4.915 0.935 ;
        RECT 6.620 1.785 6.790 1.955 ;
        RECT 6.630 0.765 6.800 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
      LAYER met1 ;
        RECT 0.580 1.940 0.870 1.985 ;
        RECT 5.145 1.940 5.435 1.985 ;
        RECT 6.560 1.940 6.850 1.985 ;
        RECT 0.580 1.800 6.850 1.940 ;
        RECT 0.580 1.755 0.870 1.800 ;
        RECT 5.145 1.755 5.435 1.800 ;
        RECT 6.560 1.755 6.850 1.800 ;
        RECT 0.990 0.920 1.280 0.965 ;
        RECT 4.685 0.920 4.975 0.965 ;
        RECT 6.570 0.920 6.860 0.965 ;
        RECT 0.990 0.780 6.860 0.920 ;
        RECT 0.990 0.735 1.280 0.780 ;
        RECT 4.685 0.735 4.975 0.780 ;
        RECT 6.570 0.735 6.860 0.780 ;
  END
END sky130_fd_sc_hd__sdfxtp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__sdfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdfxtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.040 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 2.460 1.355 2.795 1.685 ;
    END
  END D
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 3.535 1.035 4.025 1.655 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 1.780 0.785 1.950 1.685 ;
        RECT 3.085 0.785 3.255 1.115 ;
        RECT 1.780 0.615 3.255 0.785 ;
        RECT 2.475 0.305 2.650 0.615 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 11.040 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.875 0.785 6.785 1.005 ;
        RECT 8.300 0.785 10.980 1.015 ;
        RECT 0.005 0.725 4.125 0.785 ;
        RECT 5.145 0.725 10.980 0.785 ;
        RECT 0.005 0.105 10.980 0.725 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 11.230 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 11.040 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 9.285 1.675 9.615 2.395 ;
        RECT 10.135 1.675 10.465 2.395 ;
        RECT 9.285 1.505 10.955 1.675 ;
        RECT 10.655 0.905 10.955 1.505 ;
        RECT 9.285 0.735 10.955 0.905 ;
        RECT 9.285 0.305 9.615 0.735 ;
        RECT 10.135 0.305 10.465 0.735 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 11.040 2.805 ;
        RECT 0.180 1.965 0.350 2.465 ;
        RECT 0.520 2.135 0.850 2.635 ;
        RECT 0.180 1.795 0.845 1.965 ;
        RECT 0.615 0.970 0.845 1.795 ;
        RECT 0.615 0.805 0.810 0.970 ;
        RECT 0.175 0.635 0.810 0.805 ;
        RECT 1.020 0.715 1.245 2.465 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.245 0.715 ;
        RECT 1.435 2.075 1.710 2.445 ;
        RECT 1.880 2.245 2.210 2.635 ;
        RECT 2.695 2.245 3.590 2.415 ;
        RECT 1.435 1.860 3.250 2.075 ;
        RECT 1.435 0.445 1.605 1.860 ;
        RECT 2.120 1.125 2.290 1.860 ;
        RECT 3.080 1.685 3.250 1.860 ;
        RECT 3.420 1.995 3.590 2.245 ;
        RECT 3.760 2.165 3.930 2.635 ;
        RECT 4.215 2.065 4.450 2.440 ;
        RECT 4.695 2.190 5.765 2.360 ;
        RECT 4.215 1.995 4.385 2.065 ;
        RECT 3.420 1.825 4.385 1.995 ;
        RECT 3.080 1.355 3.275 1.685 ;
        RECT 2.120 0.955 2.465 1.125 ;
        RECT 4.215 0.865 4.385 1.825 ;
        RECT 3.425 0.695 4.385 0.865 ;
        RECT 4.555 1.035 4.795 1.905 ;
        RECT 4.985 1.655 5.425 2.010 ;
        RECT 5.595 1.575 5.765 2.190 ;
        RECT 5.935 1.835 6.105 2.635 ;
        RECT 6.275 2.135 6.525 2.465 ;
        RECT 6.750 2.165 7.635 2.335 ;
        RECT 5.595 1.485 6.105 1.575 ;
        RECT 5.305 1.315 6.105 1.485 ;
        RECT 4.555 0.705 5.135 1.035 ;
        RECT 3.425 0.445 3.595 0.695 ;
        RECT 4.215 0.535 4.385 0.695 ;
        RECT 5.305 0.535 5.475 1.315 ;
        RECT 5.935 1.245 6.105 1.315 ;
        RECT 5.645 1.065 5.815 1.095 ;
        RECT 6.275 1.065 6.445 2.135 ;
        RECT 6.615 1.245 6.805 1.965 ;
        RECT 6.975 1.575 7.295 1.905 ;
        RECT 5.645 0.765 6.445 1.065 ;
        RECT 6.975 1.035 7.165 1.575 ;
        RECT 7.465 1.405 7.635 2.165 ;
        RECT 7.815 2.135 8.120 2.635 ;
        RECT 8.470 1.905 8.755 2.455 ;
        RECT 7.805 1.575 8.755 1.905 ;
        RECT 8.925 1.625 9.105 2.635 ;
        RECT 9.795 1.845 9.965 2.635 ;
        RECT 10.635 1.845 10.805 2.635 ;
        RECT 1.435 0.275 1.805 0.445 ;
        RECT 1.975 0.085 2.305 0.445 ;
        RECT 2.820 0.275 3.595 0.445 ;
        RECT 3.765 0.085 3.965 0.525 ;
        RECT 4.215 0.365 4.565 0.535 ;
        RECT 4.735 0.365 5.475 0.535 ;
        RECT 5.725 0.085 6.095 0.585 ;
        RECT 6.275 0.535 6.445 0.765 ;
        RECT 6.615 0.705 7.165 1.035 ;
        RECT 7.335 1.325 7.635 1.405 ;
        RECT 8.570 1.325 8.755 1.575 ;
        RECT 7.335 0.995 8.400 1.325 ;
        RECT 8.570 1.075 10.485 1.325 ;
        RECT 7.335 0.535 7.505 0.995 ;
        RECT 8.570 0.825 8.750 1.075 ;
        RECT 6.275 0.365 6.735 0.535 ;
        RECT 6.965 0.365 7.505 0.535 ;
        RECT 7.750 0.085 8.120 0.615 ;
        RECT 8.390 0.300 8.750 0.825 ;
        RECT 8.925 0.085 9.095 0.695 ;
        RECT 9.795 0.085 9.965 0.565 ;
        RECT 10.635 0.085 10.805 0.565 ;
        RECT 0.000 -0.085 11.040 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 0.615 1.785 0.785 1.955 ;
        RECT 1.055 0.765 1.225 0.935 ;
        RECT 5.215 1.785 5.385 1.955 ;
        RECT 4.755 0.765 4.925 0.935 ;
        RECT 6.625 1.785 6.795 1.955 ;
        RECT 6.625 0.765 6.795 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
      LAYER met1 ;
        RECT 0.555 1.940 0.845 1.985 ;
        RECT 5.155 1.940 5.445 1.985 ;
        RECT 6.565 1.940 6.855 1.985 ;
        RECT 0.555 1.800 6.855 1.940 ;
        RECT 0.555 1.755 0.845 1.800 ;
        RECT 5.155 1.755 5.445 1.800 ;
        RECT 6.565 1.755 6.855 1.800 ;
        RECT 0.995 0.920 1.285 0.965 ;
        RECT 4.695 0.920 4.985 0.965 ;
        RECT 6.565 0.920 6.855 0.965 ;
        RECT 0.995 0.780 6.855 0.920 ;
        RECT 0.995 0.735 1.285 0.780 ;
        RECT 4.695 0.735 4.985 0.780 ;
        RECT 6.565 0.735 6.855 0.780 ;
  END
END sky130_fd_sc_hd__sdfxtp_4

#--------EOF---------

MACRO sky130_fd_sc_hd__sdlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdlclkp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 4.710 1.265 4.930 1.325 ;
        RECT 4.710 0.955 6.010 1.265 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.880 1.445 1.235 1.955 ;
        RECT 0.880 1.325 1.190 1.445 ;
        RECT 0.850 0.955 1.190 1.325 ;
    END
  END GATE
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.340 1.665 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.525 0.785 3.560 1.015 ;
        RECT 5.975 0.785 6.895 1.015 ;
        RECT 0.005 0.105 6.895 0.785 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 6.530 1.495 6.815 2.465 ;
        RECT 6.645 0.825 6.815 1.495 ;
        RECT 6.530 0.255 6.815 0.825 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 0.085 1.835 0.345 2.635 ;
        RECT 0.540 2.125 1.255 2.465 ;
        RECT 1.425 2.125 2.200 2.465 ;
        RECT 0.540 1.755 0.710 2.125 ;
        RECT 0.510 1.460 0.710 1.755 ;
        RECT 0.510 0.785 0.680 1.460 ;
        RECT 1.405 1.325 1.860 1.955 ;
        RECT 1.360 1.205 1.860 1.325 ;
        RECT 2.030 1.375 2.200 2.125 ;
        RECT 2.370 2.075 3.010 2.635 ;
        RECT 3.180 2.085 3.400 2.465 ;
        RECT 3.580 2.255 5.490 2.635 ;
        RECT 5.660 2.085 5.830 2.465 ;
        RECT 6.030 2.255 6.360 2.635 ;
        RECT 3.180 1.915 5.450 2.085 ;
        RECT 3.180 1.905 3.400 1.915 ;
        RECT 2.370 1.635 3.400 1.905 ;
        RECT 2.370 1.575 2.540 1.635 ;
        RECT 2.030 1.205 3.010 1.375 ;
        RECT 0.085 0.615 1.190 0.785 ;
        RECT 1.360 0.705 1.700 1.205 ;
        RECT 1.870 0.705 2.155 1.035 ;
        RECT 2.325 0.995 3.010 1.205 ;
        RECT 0.085 0.255 0.345 0.615 ;
        RECT 0.515 0.085 0.845 0.445 ;
        RECT 1.015 0.255 1.190 0.615 ;
        RECT 2.325 0.535 2.495 0.995 ;
        RECT 1.360 0.255 2.495 0.535 ;
        RECT 2.665 0.085 3.010 0.825 ;
        RECT 3.180 0.255 3.400 1.635 ;
        RECT 3.580 1.575 3.990 1.745 ;
        RECT 3.580 0.935 3.750 1.575 ;
        RECT 4.160 1.495 4.960 1.745 ;
        RECT 5.140 1.605 5.450 1.915 ;
        RECT 5.660 1.775 6.360 2.085 ;
        RECT 4.160 1.275 4.465 1.495 ;
        RECT 5.140 1.435 5.610 1.605 ;
        RECT 5.780 1.435 6.360 1.775 ;
        RECT 3.920 1.105 4.465 1.275 ;
        RECT 3.580 0.765 4.005 0.935 ;
        RECT 4.175 0.785 4.465 1.105 ;
        RECT 6.190 1.325 6.360 1.435 ;
        RECT 6.190 0.995 6.460 1.325 ;
        RECT 6.190 0.785 6.360 0.995 ;
        RECT 3.580 0.255 3.910 0.765 ;
        RECT 4.175 0.615 4.830 0.785 ;
        RECT 4.080 0.085 4.410 0.445 ;
        RECT 4.580 0.255 4.830 0.615 ;
        RECT 5.010 0.615 6.360 0.785 ;
        RECT 5.010 0.255 5.270 0.615 ;
        RECT 5.505 0.085 6.360 0.445 ;
        RECT 0.000 -0.085 6.900 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 1.525 1.445 1.695 1.615 ;
        RECT 1.985 0.765 2.155 0.935 ;
        RECT 4.295 1.445 4.465 1.615 ;
        RECT 3.835 0.765 4.005 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
      LAYER met1 ;
        RECT 1.465 1.600 1.755 1.645 ;
        RECT 4.235 1.600 4.525 1.645 ;
        RECT 1.465 1.460 4.525 1.600 ;
        RECT 1.465 1.415 1.755 1.460 ;
        RECT 4.235 1.415 4.525 1.460 ;
        RECT 1.925 0.920 2.215 0.965 ;
        RECT 3.775 0.920 4.065 0.965 ;
        RECT 1.925 0.780 4.065 0.920 ;
        RECT 1.925 0.735 2.215 0.780 ;
        RECT 3.775 0.735 4.065 0.780 ;
  END
END sky130_fd_sc_hd__sdlclkp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__sdlclkp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdlclkp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.360 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 4.705 1.265 4.925 1.325 ;
        RECT 4.705 0.955 6.050 1.265 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.855 1.445 1.240 1.955 ;
        RECT 0.855 0.955 1.195 1.445 ;
    END
  END GATE
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.340 1.665 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 7.360 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.530 0.785 3.575 1.015 ;
        RECT 6.015 0.785 7.355 1.015 ;
        RECT 0.005 0.105 7.355 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.550 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 7.360 2.960 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 6.570 1.495 6.840 2.465 ;
        RECT 6.670 1.315 6.840 1.495 ;
        RECT 6.670 1.055 7.275 1.315 ;
        RECT 6.670 0.825 6.840 1.055 ;
        RECT 6.570 0.255 6.840 0.825 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 7.360 2.805 ;
        RECT 0.085 1.835 0.345 2.635 ;
        RECT 0.515 2.125 1.260 2.465 ;
        RECT 1.430 2.125 2.205 2.465 ;
        RECT 0.515 0.785 0.685 2.125 ;
        RECT 1.410 1.325 1.865 1.955 ;
        RECT 1.365 1.205 1.865 1.325 ;
        RECT 2.035 1.375 2.205 2.125 ;
        RECT 2.375 2.075 3.015 2.635 ;
        RECT 3.185 2.085 3.405 2.465 ;
        RECT 3.575 2.255 5.530 2.635 ;
        RECT 5.700 2.085 5.870 2.465 ;
        RECT 6.070 2.255 6.400 2.635 ;
        RECT 3.185 1.915 5.490 2.085 ;
        RECT 3.185 1.905 3.405 1.915 ;
        RECT 2.375 1.635 3.405 1.905 ;
        RECT 2.375 1.575 2.545 1.635 ;
        RECT 2.035 1.205 3.015 1.375 ;
        RECT 0.085 0.615 1.195 0.785 ;
        RECT 1.365 0.705 1.705 1.205 ;
        RECT 1.875 0.705 2.160 1.035 ;
        RECT 2.330 0.995 3.015 1.205 ;
        RECT 0.085 0.255 0.345 0.615 ;
        RECT 0.515 0.085 0.845 0.445 ;
        RECT 1.015 0.255 1.195 0.615 ;
        RECT 2.330 0.535 2.500 0.995 ;
        RECT 1.365 0.255 2.500 0.535 ;
        RECT 2.670 0.085 3.015 0.825 ;
        RECT 3.185 0.255 3.405 1.635 ;
        RECT 3.575 1.575 4.040 1.745 ;
        RECT 3.575 0.935 3.745 1.575 ;
        RECT 4.210 1.495 5.010 1.745 ;
        RECT 5.180 1.605 5.490 1.915 ;
        RECT 5.700 1.775 6.400 2.085 ;
        RECT 4.210 1.275 4.460 1.495 ;
        RECT 5.180 1.435 5.650 1.605 ;
        RECT 5.820 1.435 6.400 1.775 ;
        RECT 7.010 1.485 7.275 2.635 ;
        RECT 3.915 1.105 4.460 1.275 ;
        RECT 3.575 0.765 4.000 0.935 ;
        RECT 4.170 0.785 4.460 1.105 ;
        RECT 6.230 1.325 6.400 1.435 ;
        RECT 6.230 0.995 6.500 1.325 ;
        RECT 6.230 0.785 6.400 0.995 ;
        RECT 3.575 0.255 3.925 0.765 ;
        RECT 4.170 0.615 4.825 0.785 ;
        RECT 4.095 0.085 4.425 0.445 ;
        RECT 4.595 0.255 4.825 0.615 ;
        RECT 5.100 0.615 6.400 0.785 ;
        RECT 5.100 0.255 5.310 0.615 ;
        RECT 5.490 0.085 6.400 0.445 ;
        RECT 7.010 0.085 7.275 0.885 ;
        RECT 0.000 -0.085 7.360 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 1.530 1.445 1.700 1.615 ;
        RECT 1.990 0.765 2.160 0.935 ;
        RECT 4.290 1.445 4.460 1.615 ;
        RECT 3.830 0.765 4.000 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
      LAYER met1 ;
        RECT 1.470 1.600 1.760 1.645 ;
        RECT 4.230 1.600 4.520 1.645 ;
        RECT 1.470 1.460 4.520 1.600 ;
        RECT 1.470 1.415 1.760 1.460 ;
        RECT 4.230 1.415 4.520 1.460 ;
        RECT 1.930 0.920 2.220 0.965 ;
        RECT 3.770 0.920 4.060 0.965 ;
        RECT 1.930 0.780 4.060 0.920 ;
        RECT 1.930 0.735 2.220 0.780 ;
        RECT 3.770 0.735 4.060 0.780 ;
  END
END sky130_fd_sc_hd__sdlclkp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__sdlclkp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sdlclkp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.406500 ;
    PORT
      LAYER met1 ;
        RECT 4.710 1.260 5.000 1.305 ;
        RECT 5.650 1.260 5.940 1.305 ;
        RECT 4.710 1.120 5.940 1.260 ;
        RECT 4.710 1.075 5.000 1.120 ;
        RECT 5.650 1.075 5.940 1.120 ;
    END
  END CLK
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.855 1.445 1.240 1.955 ;
        RECT 0.855 0.955 1.195 1.445 ;
    END
  END GATE
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 0.955 0.345 1.665 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 2.530 0.785 3.575 1.015 ;
        RECT 5.095 0.785 8.230 1.015 ;
        RECT 0.005 0.105 8.230 0.785 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN GCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 6.580 1.655 6.830 2.465 ;
        RECT 6.580 1.485 7.220 1.655 ;
        RECT 7.050 1.315 7.220 1.485 ;
        RECT 7.420 1.315 7.720 2.465 ;
        RECT 7.050 1.055 8.195 1.315 ;
        RECT 7.050 0.885 7.220 1.055 ;
        RECT 6.580 0.715 7.220 0.885 ;
        RECT 6.580 0.445 6.830 0.715 ;
        RECT 6.500 0.255 6.830 0.445 ;
        RECT 7.420 0.255 7.720 1.055 ;
    END
  END GCLK
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.085 1.835 0.345 2.635 ;
        RECT 0.515 2.125 1.260 2.465 ;
        RECT 1.430 2.125 2.205 2.465 ;
        RECT 0.515 0.785 0.685 2.125 ;
        RECT 1.410 1.325 1.865 1.955 ;
        RECT 1.365 1.205 1.865 1.325 ;
        RECT 2.035 1.375 2.205 2.125 ;
        RECT 2.375 2.075 3.015 2.635 ;
        RECT 3.185 2.085 3.405 2.465 ;
        RECT 3.595 2.255 5.515 2.635 ;
        RECT 5.685 2.085 5.855 2.465 ;
        RECT 6.055 2.255 6.385 2.635 ;
        RECT 3.185 1.915 5.515 2.085 ;
        RECT 3.185 1.905 3.405 1.915 ;
        RECT 2.375 1.635 3.405 1.905 ;
        RECT 2.375 1.575 2.545 1.635 ;
        RECT 2.035 1.205 3.015 1.375 ;
        RECT 0.085 0.615 1.195 0.785 ;
        RECT 1.365 0.705 1.705 1.205 ;
        RECT 1.875 0.705 2.160 1.035 ;
        RECT 2.330 0.995 3.015 1.205 ;
        RECT 0.085 0.255 0.345 0.615 ;
        RECT 0.515 0.085 0.845 0.445 ;
        RECT 1.015 0.255 1.195 0.615 ;
        RECT 2.330 0.535 2.500 0.995 ;
        RECT 1.365 0.255 2.500 0.535 ;
        RECT 2.670 0.085 3.015 0.825 ;
        RECT 3.185 0.255 3.405 1.635 ;
        RECT 3.595 1.575 4.005 1.745 ;
        RECT 3.595 0.935 3.765 1.575 ;
        RECT 4.175 1.495 4.975 1.745 ;
        RECT 4.175 1.275 4.480 1.495 ;
        RECT 3.935 1.105 4.480 1.275 ;
        RECT 3.595 0.765 4.020 0.935 ;
        RECT 4.190 0.785 4.480 1.105 ;
        RECT 4.725 0.995 4.945 1.325 ;
        RECT 5.165 0.995 5.515 1.915 ;
        RECT 5.685 1.495 6.410 2.085 ;
        RECT 7.000 1.825 7.250 2.635 ;
        RECT 5.685 0.995 6.065 1.325 ;
        RECT 6.240 1.315 6.410 1.495 ;
        RECT 7.890 1.485 8.195 2.635 ;
        RECT 6.240 1.055 6.880 1.315 ;
        RECT 6.240 0.785 6.410 1.055 ;
        RECT 3.595 0.255 3.925 0.765 ;
        RECT 4.190 0.615 4.845 0.785 ;
        RECT 4.095 0.085 4.425 0.445 ;
        RECT 4.595 0.255 4.845 0.615 ;
        RECT 5.015 0.615 6.410 0.785 ;
        RECT 5.015 0.255 5.435 0.615 ;
        RECT 5.605 0.085 6.330 0.445 ;
        RECT 7.000 0.085 7.250 0.545 ;
        RECT 7.890 0.085 8.195 0.885 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 1.530 1.445 1.700 1.615 ;
        RECT 1.990 0.765 2.160 0.935 ;
        RECT 4.310 1.445 4.480 1.615 ;
        RECT 3.850 0.765 4.020 0.935 ;
        RECT 4.770 1.105 4.940 1.275 ;
        RECT 5.710 1.105 5.880 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
      LAYER met1 ;
        RECT 1.470 1.600 1.760 1.645 ;
        RECT 4.250 1.600 4.540 1.645 ;
        RECT 1.470 1.460 4.540 1.600 ;
        RECT 1.470 1.415 1.760 1.460 ;
        RECT 4.250 1.415 4.540 1.460 ;
        RECT 1.930 0.920 2.220 0.965 ;
        RECT 3.790 0.920 4.080 0.965 ;
        RECT 1.930 0.780 4.080 0.920 ;
        RECT 1.930 0.735 2.220 0.780 ;
        RECT 3.790 0.735 4.080 0.780 ;
  END
END sky130_fd_sc_hd__sdlclkp_4

#--------EOF---------

MACRO sky130_fd_sc_hd__sedfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxbp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.260 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.720 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 2.110 1.185 2.325 1.370 ;
        RECT 2.110 0.765 2.565 1.185 ;
    END
  END DE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 5.760 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.250 1.615 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 14.260 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.170 0.785 7.135 1.145 ;
        RECT 8.400 0.785 9.320 1.005 ;
        RECT 11.305 0.785 13.955 1.015 ;
        RECT 0.005 0.465 13.955 0.785 ;
        RECT 0.005 0.105 4.965 0.465 ;
        RECT 6.435 0.105 13.955 0.465 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.435 14.450 2.910 ;
        RECT -0.190 1.305 4.885 1.435 ;
        RECT 7.200 1.305 14.450 1.435 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 14.260 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER li1 ;
        RECT 13.525 0.255 13.855 2.420 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 11.700 1.410 12.030 2.465 ;
        RECT 11.700 1.065 12.145 1.410 ;
        RECT 11.815 0.255 12.145 1.065 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 14.260 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.845 1.965 ;
        RECT 0.615 0.805 0.845 1.795 ;
        RECT 0.175 0.635 0.845 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 2.465 ;
        RECT 1.355 1.890 1.785 2.465 ;
        RECT 2.235 1.890 2.565 2.635 ;
        RECT 1.355 0.515 1.525 1.890 ;
        RECT 2.755 1.720 3.085 2.425 ;
        RECT 3.265 1.825 3.460 2.635 ;
        RECT 4.125 2.020 4.455 2.465 ;
        RECT 4.635 2.210 4.965 2.465 ;
        RECT 4.125 1.820 4.515 2.020 ;
        RECT 2.495 1.355 3.085 1.720 ;
        RECT 2.780 1.175 3.085 1.355 ;
        RECT 3.805 1.320 4.175 1.650 ;
        RECT 2.780 0.845 3.635 1.175 ;
        RECT 1.355 0.255 1.785 0.515 ;
        RECT 2.235 0.085 2.565 0.515 ;
        RECT 2.780 0.255 3.005 0.845 ;
        RECT 3.805 0.685 3.975 1.320 ;
        RECT 4.345 1.150 4.515 1.820 ;
        RECT 4.145 0.980 4.515 1.150 ;
        RECT 4.685 1.785 4.965 2.210 ;
        RECT 5.155 2.005 5.495 2.465 ;
        RECT 5.665 2.175 6.010 2.635 ;
        RECT 6.675 2.150 7.005 2.465 ;
        RECT 7.215 2.175 8.255 2.375 ;
        RECT 5.155 1.835 6.585 2.005 ;
        RECT 3.185 0.085 3.515 0.610 ;
        RECT 4.145 0.255 4.415 0.980 ;
        RECT 4.685 0.825 4.855 1.785 ;
        RECT 5.420 0.935 5.590 1.835 ;
        RECT 6.385 1.355 6.585 1.835 ;
        RECT 6.755 1.865 7.005 2.150 ;
        RECT 6.755 1.185 6.925 1.865 ;
        RECT 4.595 0.645 4.855 0.825 ;
        RECT 4.595 0.255 4.795 0.645 ;
        RECT 5.260 0.515 5.590 0.935 ;
        RECT 4.965 0.255 5.590 0.515 ;
        RECT 5.760 0.085 6.010 0.905 ;
        RECT 6.515 0.565 6.925 1.185 ;
        RECT 7.095 1.125 7.280 1.720 ;
        RECT 7.450 1.655 7.915 2.005 ;
        RECT 7.450 0.955 7.620 1.655 ;
        RECT 8.085 1.575 8.255 2.175 ;
        RECT 8.425 1.835 8.660 2.635 ;
        RECT 8.085 1.485 8.660 1.575 ;
        RECT 7.115 0.735 7.620 0.955 ;
        RECT 7.810 1.315 8.660 1.485 ;
        RECT 7.810 0.565 7.980 1.315 ;
        RECT 8.490 1.245 8.660 1.315 ;
        RECT 8.830 1.375 9.160 2.465 ;
        RECT 9.370 2.105 9.660 2.635 ;
        RECT 10.225 2.165 11.190 2.355 ;
        RECT 8.170 1.065 8.370 1.095 ;
        RECT 8.830 1.065 9.745 1.375 ;
        RECT 10.090 1.245 10.280 1.965 ;
        RECT 8.170 1.045 9.745 1.065 ;
        RECT 8.170 0.765 9.235 1.045 ;
        RECT 10.450 1.035 10.770 1.995 ;
        RECT 6.515 0.255 7.135 0.565 ;
        RECT 7.305 0.255 7.980 0.565 ;
        RECT 8.245 0.085 8.640 0.560 ;
        RECT 8.830 0.255 9.235 0.765 ;
        RECT 10.305 0.705 10.770 1.035 ;
        RECT 9.465 0.085 9.740 0.615 ;
        RECT 10.940 0.535 11.190 2.165 ;
        RECT 11.360 1.495 11.530 2.635 ;
        RECT 12.200 1.575 12.430 2.010 ;
        RECT 12.600 1.220 12.940 2.465 ;
        RECT 13.110 1.465 13.355 2.635 ;
        RECT 10.325 0.330 11.190 0.535 ;
        RECT 11.395 0.085 11.645 0.900 ;
        RECT 12.315 0.890 12.940 1.220 ;
        RECT 12.600 0.255 12.940 0.890 ;
        RECT 13.110 0.085 13.355 0.900 ;
        RECT 0.000 -0.085 14.260 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 0.635 1.785 0.805 1.955 ;
        RECT 1.015 1.445 1.185 1.615 ;
        RECT 1.355 0.425 1.525 0.595 ;
        RECT 3.805 0.765 3.975 0.935 ;
        RECT 7.510 1.785 7.680 1.955 ;
        RECT 4.185 0.425 4.355 0.595 ;
        RECT 4.615 0.425 4.785 0.595 ;
        RECT 7.100 1.445 7.270 1.615 ;
        RECT 6.530 0.425 6.700 0.595 ;
        RECT 10.100 1.785 10.270 1.955 ;
        RECT 10.520 1.445 10.690 1.615 ;
        RECT 10.980 1.785 11.150 1.955 ;
        RECT 12.230 1.785 12.400 1.955 ;
        RECT 12.690 0.765 12.860 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
      LAYER met1 ;
        RECT 0.575 1.940 0.865 1.985 ;
        RECT 7.450 1.940 7.740 1.985 ;
        RECT 10.040 1.940 10.330 1.985 ;
        RECT 0.575 1.800 10.330 1.940 ;
        RECT 0.575 1.755 0.865 1.800 ;
        RECT 7.450 1.755 7.740 1.800 ;
        RECT 10.040 1.755 10.330 1.800 ;
        RECT 10.920 1.940 11.210 1.985 ;
        RECT 12.170 1.940 12.460 1.985 ;
        RECT 10.920 1.800 12.460 1.940 ;
        RECT 10.920 1.755 11.210 1.800 ;
        RECT 12.170 1.755 12.460 1.800 ;
        RECT 0.955 1.600 1.245 1.645 ;
        RECT 7.040 1.600 7.330 1.645 ;
        RECT 10.460 1.600 10.750 1.645 ;
        RECT 0.955 1.460 10.750 1.600 ;
        RECT 0.955 1.415 1.245 1.460 ;
        RECT 7.040 1.415 7.330 1.460 ;
        RECT 10.460 1.415 10.750 1.460 ;
        RECT 3.745 0.920 4.035 0.965 ;
        RECT 12.630 0.920 12.920 0.965 ;
        RECT 3.745 0.780 12.920 0.920 ;
        RECT 3.745 0.735 4.035 0.780 ;
        RECT 12.630 0.735 12.920 0.780 ;
        RECT 1.295 0.580 1.585 0.625 ;
        RECT 4.125 0.580 4.415 0.625 ;
        RECT 1.295 0.395 4.415 0.580 ;
        RECT 4.555 0.580 4.845 0.625 ;
        RECT 6.470 0.580 6.760 0.625 ;
        RECT 4.555 0.395 6.760 0.580 ;
  END
END sky130_fd_sc_hd__sedfxbp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__sedfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxbp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.180 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.720 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 2.110 1.185 2.325 1.370 ;
        RECT 2.110 0.765 2.565 1.185 ;
    END
  END DE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 5.760 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.250 1.615 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 15.180 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.170 0.785 7.135 1.145 ;
        RECT 8.400 0.785 9.320 1.005 ;
        RECT 11.305 0.785 14.795 1.015 ;
        RECT 0.005 0.465 14.795 0.785 ;
        RECT 0.005 0.105 4.965 0.465 ;
        RECT 6.435 0.105 14.795 0.465 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.435 15.370 2.910 ;
        RECT -0.190 1.305 4.885 1.435 ;
        RECT 7.200 1.305 15.370 1.435 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 15.180 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 13.935 0.255 14.265 2.420 ;
    END
  END Q
  PIN Q_N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 11.700 1.300 12.030 2.465 ;
        RECT 11.700 1.065 12.145 1.300 ;
        RECT 11.815 0.255 12.145 1.065 ;
    END
  END Q_N
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 15.180 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.845 1.965 ;
        RECT 0.615 0.805 0.845 1.795 ;
        RECT 0.175 0.635 0.845 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 2.465 ;
        RECT 1.355 1.890 1.785 2.465 ;
        RECT 2.235 1.890 2.565 2.635 ;
        RECT 1.355 0.515 1.525 1.890 ;
        RECT 2.755 1.720 3.085 2.425 ;
        RECT 3.265 1.825 3.460 2.635 ;
        RECT 4.125 2.020 4.455 2.465 ;
        RECT 4.635 2.210 4.965 2.465 ;
        RECT 4.125 1.820 4.515 2.020 ;
        RECT 2.495 1.355 3.085 1.720 ;
        RECT 2.780 1.175 3.085 1.355 ;
        RECT 3.805 1.320 4.175 1.650 ;
        RECT 2.780 0.845 3.635 1.175 ;
        RECT 1.355 0.255 1.785 0.515 ;
        RECT 2.235 0.085 2.565 0.515 ;
        RECT 2.780 0.255 3.005 0.845 ;
        RECT 3.805 0.685 3.975 1.320 ;
        RECT 4.345 1.150 4.515 1.820 ;
        RECT 4.145 0.980 4.515 1.150 ;
        RECT 4.685 1.785 4.965 2.210 ;
        RECT 5.155 2.005 5.495 2.465 ;
        RECT 5.665 2.175 6.010 2.635 ;
        RECT 6.675 2.150 7.005 2.465 ;
        RECT 7.215 2.175 8.255 2.375 ;
        RECT 5.155 1.835 6.585 2.005 ;
        RECT 3.185 0.085 3.515 0.610 ;
        RECT 4.145 0.255 4.415 0.980 ;
        RECT 4.685 0.825 4.855 1.785 ;
        RECT 5.420 0.935 5.590 1.835 ;
        RECT 6.385 1.355 6.585 1.835 ;
        RECT 6.755 1.865 7.005 2.150 ;
        RECT 6.755 1.185 6.925 1.865 ;
        RECT 4.595 0.645 4.855 0.825 ;
        RECT 4.595 0.255 4.795 0.645 ;
        RECT 5.260 0.515 5.590 0.935 ;
        RECT 4.965 0.255 5.590 0.515 ;
        RECT 5.760 0.085 6.010 0.905 ;
        RECT 6.515 0.565 6.925 1.185 ;
        RECT 7.095 1.125 7.280 1.720 ;
        RECT 7.450 1.655 7.915 2.005 ;
        RECT 7.450 0.955 7.620 1.655 ;
        RECT 8.085 1.575 8.255 2.175 ;
        RECT 8.425 1.835 8.660 2.635 ;
        RECT 8.085 1.485 8.660 1.575 ;
        RECT 7.115 0.735 7.620 0.955 ;
        RECT 7.810 1.315 8.660 1.485 ;
        RECT 7.810 0.565 7.980 1.315 ;
        RECT 8.490 1.245 8.660 1.315 ;
        RECT 8.830 1.375 9.160 2.465 ;
        RECT 9.370 2.105 9.660 2.635 ;
        RECT 10.225 2.165 11.190 2.355 ;
        RECT 8.170 1.065 8.370 1.095 ;
        RECT 8.830 1.065 9.745 1.375 ;
        RECT 10.090 1.245 10.280 1.965 ;
        RECT 8.170 1.045 9.745 1.065 ;
        RECT 8.170 0.765 9.235 1.045 ;
        RECT 10.450 1.035 10.770 1.995 ;
        RECT 6.515 0.255 7.135 0.565 ;
        RECT 7.305 0.255 7.980 0.565 ;
        RECT 8.245 0.085 8.640 0.560 ;
        RECT 8.830 0.255 9.235 0.765 ;
        RECT 10.305 0.705 10.770 1.035 ;
        RECT 9.465 0.085 9.740 0.615 ;
        RECT 10.940 0.535 11.190 2.165 ;
        RECT 11.360 1.495 11.530 2.635 ;
        RECT 12.200 1.465 12.450 2.635 ;
        RECT 12.620 1.575 12.850 2.010 ;
        RECT 13.020 1.220 13.360 2.465 ;
        RECT 13.530 1.465 13.765 2.635 ;
        RECT 14.435 1.465 14.695 2.635 ;
        RECT 10.325 0.330 11.190 0.535 ;
        RECT 11.395 0.085 11.645 0.900 ;
        RECT 12.315 0.085 12.565 0.900 ;
        RECT 12.735 0.890 13.360 1.220 ;
        RECT 13.020 0.255 13.360 0.890 ;
        RECT 13.530 0.085 13.765 0.900 ;
        RECT 14.435 0.085 14.695 0.900 ;
        RECT 0.000 -0.085 15.180 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 14.865 2.635 15.035 2.805 ;
        RECT 0.635 1.785 0.805 1.955 ;
        RECT 1.015 1.445 1.185 1.615 ;
        RECT 1.355 0.425 1.525 0.595 ;
        RECT 3.805 0.765 3.975 0.935 ;
        RECT 7.510 1.785 7.680 1.955 ;
        RECT 4.185 0.425 4.355 0.595 ;
        RECT 4.615 0.425 4.785 0.595 ;
        RECT 7.100 1.445 7.270 1.615 ;
        RECT 6.530 0.425 6.700 0.595 ;
        RECT 10.100 1.785 10.270 1.955 ;
        RECT 10.520 1.445 10.690 1.615 ;
        RECT 10.980 1.785 11.150 1.955 ;
        RECT 12.650 1.785 12.820 1.955 ;
        RECT 13.110 0.765 13.280 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
        RECT 14.865 -0.085 15.035 0.085 ;
      LAYER met1 ;
        RECT 0.575 1.940 0.865 1.985 ;
        RECT 7.450 1.940 7.740 1.985 ;
        RECT 10.040 1.940 10.330 1.985 ;
        RECT 0.575 1.800 10.330 1.940 ;
        RECT 0.575 1.755 0.865 1.800 ;
        RECT 7.450 1.755 7.740 1.800 ;
        RECT 10.040 1.755 10.330 1.800 ;
        RECT 10.920 1.940 11.210 1.985 ;
        RECT 12.590 1.940 12.880 1.985 ;
        RECT 10.920 1.800 12.880 1.940 ;
        RECT 10.920 1.755 11.210 1.800 ;
        RECT 12.590 1.755 12.880 1.800 ;
        RECT 0.955 1.600 1.245 1.645 ;
        RECT 7.040 1.600 7.330 1.645 ;
        RECT 10.460 1.600 10.750 1.645 ;
        RECT 0.955 1.460 10.750 1.600 ;
        RECT 0.955 1.415 1.245 1.460 ;
        RECT 7.040 1.415 7.330 1.460 ;
        RECT 10.460 1.415 10.750 1.460 ;
        RECT 3.745 0.920 4.035 0.965 ;
        RECT 13.050 0.920 13.340 0.965 ;
        RECT 3.745 0.780 13.340 0.920 ;
        RECT 3.745 0.735 4.035 0.780 ;
        RECT 13.050 0.735 13.340 0.780 ;
        RECT 1.295 0.580 1.585 0.625 ;
        RECT 4.125 0.580 4.415 0.625 ;
        RECT 1.295 0.395 4.415 0.580 ;
        RECT 4.555 0.580 4.845 0.625 ;
        RECT 6.470 0.580 6.760 0.625 ;
        RECT 4.555 0.395 6.760 0.580 ;
  END
END sky130_fd_sc_hd__sedfxbp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__sedfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.340 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.720 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 2.110 1.185 2.325 1.370 ;
        RECT 2.110 0.765 2.565 1.185 ;
    END
  END DE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 5.760 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.250 1.615 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 13.340 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.170 0.785 7.135 1.145 ;
        RECT 8.400 0.785 9.320 1.005 ;
        RECT 12.245 0.785 13.195 1.015 ;
        RECT 0.005 0.465 13.195 0.785 ;
        RECT 0.005 0.105 4.965 0.465 ;
        RECT 6.435 0.105 13.195 0.465 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.435 13.530 2.910 ;
        RECT -0.190 1.305 4.885 1.435 ;
        RECT 7.200 1.305 13.530 1.435 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 13.340 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.462000 ;
    PORT
      LAYER li1 ;
        RECT 12.765 0.305 13.095 2.420 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 13.340 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.845 1.965 ;
        RECT 0.615 0.805 0.845 1.795 ;
        RECT 0.175 0.635 0.845 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 2.465 ;
        RECT 1.355 1.890 1.785 2.465 ;
        RECT 2.235 1.890 2.565 2.635 ;
        RECT 1.355 0.515 1.525 1.890 ;
        RECT 2.755 1.720 3.085 2.425 ;
        RECT 3.265 1.825 3.460 2.635 ;
        RECT 4.125 2.020 4.455 2.465 ;
        RECT 4.635 2.210 4.965 2.465 ;
        RECT 4.125 1.820 4.515 2.020 ;
        RECT 2.495 1.355 3.085 1.720 ;
        RECT 2.780 1.175 3.085 1.355 ;
        RECT 3.805 1.320 4.175 1.650 ;
        RECT 2.780 0.845 3.635 1.175 ;
        RECT 1.355 0.255 1.785 0.515 ;
        RECT 2.235 0.085 2.565 0.515 ;
        RECT 2.780 0.255 3.005 0.845 ;
        RECT 3.805 0.685 3.975 1.320 ;
        RECT 4.345 1.150 4.515 1.820 ;
        RECT 4.145 0.980 4.515 1.150 ;
        RECT 4.685 1.785 4.965 2.210 ;
        RECT 5.155 2.005 5.495 2.465 ;
        RECT 5.665 2.175 6.010 2.635 ;
        RECT 6.675 2.150 7.005 2.465 ;
        RECT 7.215 2.175 8.255 2.375 ;
        RECT 5.155 1.835 6.585 2.005 ;
        RECT 3.185 0.085 3.515 0.610 ;
        RECT 4.145 0.255 4.415 0.980 ;
        RECT 4.685 0.825 4.855 1.785 ;
        RECT 5.420 0.935 5.590 1.835 ;
        RECT 6.385 1.355 6.585 1.835 ;
        RECT 6.755 1.865 7.005 2.150 ;
        RECT 6.755 1.185 6.925 1.865 ;
        RECT 4.595 0.645 4.855 0.825 ;
        RECT 4.595 0.255 4.795 0.645 ;
        RECT 5.260 0.515 5.590 0.935 ;
        RECT 4.965 0.255 5.590 0.515 ;
        RECT 5.760 0.085 6.010 0.905 ;
        RECT 6.515 0.565 6.925 1.185 ;
        RECT 7.095 1.125 7.280 1.720 ;
        RECT 7.450 1.655 7.915 2.005 ;
        RECT 7.450 0.955 7.620 1.655 ;
        RECT 8.085 1.575 8.255 2.175 ;
        RECT 8.425 1.835 8.660 2.635 ;
        RECT 8.085 1.485 8.660 1.575 ;
        RECT 7.115 0.735 7.620 0.955 ;
        RECT 7.810 1.315 8.660 1.485 ;
        RECT 7.810 0.565 7.980 1.315 ;
        RECT 8.490 1.245 8.660 1.315 ;
        RECT 8.830 1.375 9.160 2.465 ;
        RECT 9.370 2.105 9.660 2.635 ;
        RECT 10.225 2.165 11.110 2.355 ;
        RECT 8.170 1.065 8.370 1.095 ;
        RECT 8.830 1.065 9.745 1.375 ;
        RECT 10.090 1.245 10.280 1.965 ;
        RECT 8.170 1.045 9.745 1.065 ;
        RECT 8.170 0.765 9.235 1.045 ;
        RECT 10.450 1.035 10.770 1.995 ;
        RECT 6.515 0.255 7.135 0.565 ;
        RECT 7.305 0.255 7.980 0.565 ;
        RECT 8.245 0.085 8.640 0.560 ;
        RECT 8.830 0.255 9.235 0.765 ;
        RECT 10.305 0.705 10.770 1.035 ;
        RECT 10.940 1.325 11.110 2.165 ;
        RECT 11.280 2.135 11.540 2.635 ;
        RECT 11.840 1.905 12.180 2.465 ;
        RECT 11.280 1.530 12.180 1.905 ;
        RECT 10.940 0.995 11.810 1.325 ;
        RECT 9.465 0.085 9.740 0.615 ;
        RECT 10.940 0.535 11.110 0.995 ;
        RECT 11.990 0.825 12.180 1.530 ;
        RECT 12.350 1.465 12.595 2.635 ;
        RECT 10.325 0.330 11.110 0.535 ;
        RECT 11.350 0.085 11.665 0.615 ;
        RECT 11.850 0.300 12.180 0.825 ;
        RECT 12.350 0.085 12.595 0.900 ;
        RECT 0.000 -0.085 13.340 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 0.635 1.785 0.805 1.955 ;
        RECT 1.015 1.445 1.185 1.615 ;
        RECT 1.355 0.425 1.525 0.595 ;
        RECT 3.805 0.765 3.975 0.935 ;
        RECT 7.510 1.785 7.680 1.955 ;
        RECT 4.185 0.425 4.355 0.595 ;
        RECT 4.615 0.425 4.785 0.595 ;
        RECT 7.100 1.445 7.270 1.615 ;
        RECT 6.530 0.425 6.700 0.595 ;
        RECT 10.100 1.785 10.270 1.955 ;
        RECT 10.520 1.445 10.690 1.615 ;
        RECT 12.000 0.765 12.170 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
      LAYER met1 ;
        RECT 0.575 1.940 0.865 1.985 ;
        RECT 7.450 1.940 7.740 1.985 ;
        RECT 10.040 1.940 10.330 1.985 ;
        RECT 0.575 1.800 10.330 1.940 ;
        RECT 0.575 1.755 0.865 1.800 ;
        RECT 7.450 1.755 7.740 1.800 ;
        RECT 10.040 1.755 10.330 1.800 ;
        RECT 0.955 1.600 1.245 1.645 ;
        RECT 7.040 1.600 7.330 1.645 ;
        RECT 10.460 1.600 10.750 1.645 ;
        RECT 0.955 1.460 10.750 1.600 ;
        RECT 0.955 1.415 1.245 1.460 ;
        RECT 7.040 1.415 7.330 1.460 ;
        RECT 10.460 1.415 10.750 1.460 ;
        RECT 3.745 0.920 4.035 0.965 ;
        RECT 11.940 0.920 12.230 0.965 ;
        RECT 3.745 0.780 12.230 0.920 ;
        RECT 3.745 0.735 4.035 0.780 ;
        RECT 11.940 0.735 12.230 0.780 ;
        RECT 1.295 0.580 1.585 0.625 ;
        RECT 4.125 0.580 4.415 0.625 ;
        RECT 1.295 0.395 4.415 0.580 ;
        RECT 4.555 0.580 4.845 0.625 ;
        RECT 6.470 0.580 6.760 0.625 ;
        RECT 4.555 0.395 6.760 0.580 ;
  END
END sky130_fd_sc_hd__sedfxtp_1

#--------EOF---------

MACRO sky130_fd_sc_hd__sedfxtp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxtp_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 13.800 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.720 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 2.110 1.185 2.325 1.370 ;
        RECT 2.110 0.765 2.565 1.185 ;
    END
  END DE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 5.760 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.250 1.615 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 13.800 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.170 0.785 7.135 1.145 ;
        RECT 8.400 0.785 9.320 1.005 ;
        RECT 12.245 0.785 13.625 1.015 ;
        RECT 0.005 0.465 13.625 0.785 ;
        RECT 0.005 0.105 4.965 0.465 ;
        RECT 6.435 0.105 13.625 0.465 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.435 13.990 2.910 ;
        RECT -0.190 1.305 4.885 1.435 ;
        RECT 7.200 1.305 13.990 1.435 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 13.800 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 12.755 0.305 13.085 2.420 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 13.800 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.845 1.965 ;
        RECT 0.615 0.805 0.845 1.795 ;
        RECT 0.175 0.635 0.845 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 2.465 ;
        RECT 1.355 1.890 1.785 2.465 ;
        RECT 2.235 1.890 2.565 2.635 ;
        RECT 1.355 0.515 1.525 1.890 ;
        RECT 2.755 1.720 3.085 2.425 ;
        RECT 3.265 1.825 3.460 2.635 ;
        RECT 4.125 2.020 4.455 2.465 ;
        RECT 4.635 2.210 4.965 2.465 ;
        RECT 4.125 1.820 4.515 2.020 ;
        RECT 2.495 1.355 3.085 1.720 ;
        RECT 2.780 1.175 3.085 1.355 ;
        RECT 3.805 1.320 4.175 1.650 ;
        RECT 2.780 0.845 3.635 1.175 ;
        RECT 1.355 0.255 1.785 0.515 ;
        RECT 2.235 0.085 2.565 0.515 ;
        RECT 2.780 0.255 3.005 0.845 ;
        RECT 3.805 0.685 3.975 1.320 ;
        RECT 4.345 1.150 4.515 1.820 ;
        RECT 4.145 0.980 4.515 1.150 ;
        RECT 4.685 1.785 4.965 2.210 ;
        RECT 5.155 2.005 5.495 2.465 ;
        RECT 5.665 2.175 6.010 2.635 ;
        RECT 6.675 2.150 7.005 2.465 ;
        RECT 7.215 2.175 8.255 2.375 ;
        RECT 5.155 1.835 6.585 2.005 ;
        RECT 3.185 0.085 3.515 0.610 ;
        RECT 4.145 0.255 4.415 0.980 ;
        RECT 4.685 0.825 4.855 1.785 ;
        RECT 5.420 0.935 5.590 1.835 ;
        RECT 6.385 1.355 6.585 1.835 ;
        RECT 6.755 1.865 7.005 2.150 ;
        RECT 6.755 1.185 6.925 1.865 ;
        RECT 4.595 0.645 4.855 0.825 ;
        RECT 4.595 0.255 4.795 0.645 ;
        RECT 5.260 0.515 5.590 0.935 ;
        RECT 4.965 0.255 5.590 0.515 ;
        RECT 5.760 0.085 6.010 0.905 ;
        RECT 6.515 0.565 6.925 1.185 ;
        RECT 7.095 1.125 7.280 1.720 ;
        RECT 7.450 1.655 7.915 2.005 ;
        RECT 7.450 0.955 7.620 1.655 ;
        RECT 8.085 1.575 8.255 2.175 ;
        RECT 8.425 1.835 8.660 2.635 ;
        RECT 8.085 1.485 8.660 1.575 ;
        RECT 7.115 0.735 7.620 0.955 ;
        RECT 7.810 1.315 8.660 1.485 ;
        RECT 7.810 0.565 7.980 1.315 ;
        RECT 8.490 1.245 8.660 1.315 ;
        RECT 8.830 1.375 9.160 2.465 ;
        RECT 9.370 2.105 9.660 2.635 ;
        RECT 10.225 2.165 11.110 2.355 ;
        RECT 8.170 1.065 8.370 1.095 ;
        RECT 8.830 1.065 9.745 1.375 ;
        RECT 10.090 1.245 10.280 1.965 ;
        RECT 8.170 1.045 9.745 1.065 ;
        RECT 8.170 0.765 9.235 1.045 ;
        RECT 10.450 1.035 10.770 1.995 ;
        RECT 6.515 0.255 7.135 0.565 ;
        RECT 7.305 0.255 7.980 0.565 ;
        RECT 8.245 0.085 8.640 0.560 ;
        RECT 8.830 0.255 9.235 0.765 ;
        RECT 10.305 0.705 10.770 1.035 ;
        RECT 10.940 1.325 11.110 2.165 ;
        RECT 11.280 2.135 11.540 2.635 ;
        RECT 11.840 1.905 12.180 2.465 ;
        RECT 11.280 1.530 12.180 1.905 ;
        RECT 10.940 0.995 11.810 1.325 ;
        RECT 9.465 0.085 9.740 0.615 ;
        RECT 10.940 0.535 11.110 0.995 ;
        RECT 11.990 0.825 12.180 1.530 ;
        RECT 12.350 1.465 12.585 2.635 ;
        RECT 13.255 1.465 13.515 2.635 ;
        RECT 10.325 0.330 11.110 0.535 ;
        RECT 11.350 0.085 11.665 0.615 ;
        RECT 11.850 0.300 12.180 0.825 ;
        RECT 12.350 0.085 12.585 0.900 ;
        RECT 13.255 0.085 13.515 0.900 ;
        RECT 0.000 -0.085 13.800 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 0.635 1.785 0.805 1.955 ;
        RECT 1.015 1.445 1.185 1.615 ;
        RECT 1.355 0.425 1.525 0.595 ;
        RECT 3.805 0.765 3.975 0.935 ;
        RECT 7.510 1.785 7.680 1.955 ;
        RECT 4.185 0.425 4.355 0.595 ;
        RECT 4.615 0.425 4.785 0.595 ;
        RECT 7.100 1.445 7.270 1.615 ;
        RECT 6.530 0.425 6.700 0.595 ;
        RECT 10.100 1.785 10.270 1.955 ;
        RECT 10.520 1.445 10.690 1.615 ;
        RECT 12.000 0.765 12.170 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
      LAYER met1 ;
        RECT 0.575 1.940 0.865 1.985 ;
        RECT 7.450 1.940 7.740 1.985 ;
        RECT 10.040 1.940 10.330 1.985 ;
        RECT 0.575 1.800 10.330 1.940 ;
        RECT 0.575 1.755 0.865 1.800 ;
        RECT 7.450 1.755 7.740 1.800 ;
        RECT 10.040 1.755 10.330 1.800 ;
        RECT 0.955 1.600 1.245 1.645 ;
        RECT 7.040 1.600 7.330 1.645 ;
        RECT 10.460 1.600 10.750 1.645 ;
        RECT 0.955 1.460 10.750 1.600 ;
        RECT 0.955 1.415 1.245 1.460 ;
        RECT 7.040 1.415 7.330 1.460 ;
        RECT 10.460 1.415 10.750 1.460 ;
        RECT 3.745 0.920 4.035 0.965 ;
        RECT 11.940 0.920 12.230 0.965 ;
        RECT 3.745 0.780 12.230 0.920 ;
        RECT 3.745 0.735 4.035 0.780 ;
        RECT 11.940 0.735 12.230 0.780 ;
        RECT 1.295 0.580 1.585 0.625 ;
        RECT 4.125 0.580 4.415 0.625 ;
        RECT 1.295 0.395 4.415 0.580 ;
        RECT 4.555 0.580 4.845 0.625 ;
        RECT 6.470 0.580 6.760 0.625 ;
        RECT 4.555 0.395 6.760 0.580 ;
  END
END sky130_fd_sc_hd__sedfxtp_2

#--------EOF---------

MACRO sky130_fd_sc_hd__sedfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__sedfxtp_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.720 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 0.095 0.975 0.445 1.625 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.695 0.765 1.915 1.720 ;
    END
  END D
  PIN DE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 2.110 1.185 2.325 1.370 ;
        RECT 2.110 0.765 2.565 1.185 ;
    END
  END DE
  PIN SCD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 5.760 1.105 6.215 1.665 ;
    END
  END SCD
  PIN SCE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.318000 ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.105 5.250 1.615 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 14.720 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 5.170 0.785 7.135 1.145 ;
        RECT 8.400 0.785 9.320 1.005 ;
        RECT 12.245 0.785 14.465 1.015 ;
        RECT 0.005 0.465 14.465 0.785 ;
        RECT 0.005 0.105 4.965 0.465 ;
        RECT 6.435 0.105 14.465 0.465 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.435 14.910 2.910 ;
        RECT -0.190 1.305 4.885 1.435 ;
        RECT 7.200 1.305 14.910 1.435 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 14.720 2.960 ;
    END
  END VPWR
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 12.755 1.295 13.085 2.420 ;
        RECT 13.595 1.295 13.925 2.420 ;
        RECT 12.755 1.070 13.925 1.295 ;
        RECT 12.755 0.305 13.085 1.070 ;
        RECT 13.595 0.305 13.925 1.070 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 14.720 2.805 ;
        RECT 0.175 1.965 0.345 2.465 ;
        RECT 0.515 2.135 0.845 2.635 ;
        RECT 0.175 1.795 0.845 1.965 ;
        RECT 0.615 0.805 0.845 1.795 ;
        RECT 0.175 0.635 0.845 0.805 ;
        RECT 0.175 0.345 0.345 0.635 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.015 0.345 1.185 2.465 ;
        RECT 1.355 1.890 1.785 2.465 ;
        RECT 2.235 1.890 2.565 2.635 ;
        RECT 1.355 0.515 1.525 1.890 ;
        RECT 2.755 1.720 3.085 2.425 ;
        RECT 3.265 1.825 3.460 2.635 ;
        RECT 4.125 2.020 4.455 2.465 ;
        RECT 4.635 2.210 4.965 2.465 ;
        RECT 4.125 1.820 4.515 2.020 ;
        RECT 2.495 1.355 3.085 1.720 ;
        RECT 2.780 1.175 3.085 1.355 ;
        RECT 3.805 1.320 4.175 1.650 ;
        RECT 2.780 0.845 3.635 1.175 ;
        RECT 1.355 0.255 1.785 0.515 ;
        RECT 2.235 0.085 2.565 0.515 ;
        RECT 2.780 0.255 3.005 0.845 ;
        RECT 3.805 0.685 3.975 1.320 ;
        RECT 4.345 1.150 4.515 1.820 ;
        RECT 4.145 0.980 4.515 1.150 ;
        RECT 4.685 1.785 4.965 2.210 ;
        RECT 5.155 2.005 5.495 2.465 ;
        RECT 5.665 2.175 6.010 2.635 ;
        RECT 6.675 2.150 7.005 2.465 ;
        RECT 7.215 2.175 8.255 2.375 ;
        RECT 5.155 1.835 6.585 2.005 ;
        RECT 3.185 0.085 3.515 0.610 ;
        RECT 4.145 0.255 4.415 0.980 ;
        RECT 4.685 0.825 4.855 1.785 ;
        RECT 5.420 0.935 5.590 1.835 ;
        RECT 6.385 1.355 6.585 1.835 ;
        RECT 6.755 1.865 7.005 2.150 ;
        RECT 6.755 1.185 6.925 1.865 ;
        RECT 4.595 0.645 4.855 0.825 ;
        RECT 4.595 0.255 4.795 0.645 ;
        RECT 5.260 0.515 5.590 0.935 ;
        RECT 4.965 0.255 5.590 0.515 ;
        RECT 5.760 0.085 6.010 0.905 ;
        RECT 6.515 0.565 6.925 1.185 ;
        RECT 7.095 1.125 7.280 1.720 ;
        RECT 7.450 1.655 7.915 2.005 ;
        RECT 7.450 0.955 7.620 1.655 ;
        RECT 8.085 1.575 8.255 2.175 ;
        RECT 8.425 1.835 8.660 2.635 ;
        RECT 8.085 1.485 8.660 1.575 ;
        RECT 7.115 0.735 7.620 0.955 ;
        RECT 7.810 1.315 8.660 1.485 ;
        RECT 7.810 0.565 7.980 1.315 ;
        RECT 8.490 1.245 8.660 1.315 ;
        RECT 8.830 1.375 9.160 2.465 ;
        RECT 9.370 2.105 9.660 2.635 ;
        RECT 10.225 2.165 11.110 2.355 ;
        RECT 8.170 1.065 8.370 1.095 ;
        RECT 8.830 1.065 9.745 1.375 ;
        RECT 10.090 1.245 10.280 1.965 ;
        RECT 8.170 1.045 9.745 1.065 ;
        RECT 8.170 0.765 9.235 1.045 ;
        RECT 10.450 1.035 10.770 1.995 ;
        RECT 6.515 0.255 7.135 0.565 ;
        RECT 7.305 0.255 7.980 0.565 ;
        RECT 8.245 0.085 8.640 0.560 ;
        RECT 8.830 0.255 9.235 0.765 ;
        RECT 10.305 0.705 10.770 1.035 ;
        RECT 10.940 1.325 11.110 2.165 ;
        RECT 11.280 2.135 11.540 2.635 ;
        RECT 11.840 1.905 12.180 2.465 ;
        RECT 11.280 1.530 12.180 1.905 ;
        RECT 10.940 0.995 11.810 1.325 ;
        RECT 9.465 0.085 9.740 0.615 ;
        RECT 10.940 0.535 11.110 0.995 ;
        RECT 11.990 0.825 12.180 1.530 ;
        RECT 12.350 1.465 12.585 2.635 ;
        RECT 13.255 1.465 13.425 2.635 ;
        RECT 14.095 1.465 14.355 2.635 ;
        RECT 10.325 0.330 11.110 0.535 ;
        RECT 11.350 0.085 11.665 0.615 ;
        RECT 11.850 0.300 12.180 0.825 ;
        RECT 12.350 0.085 12.585 0.900 ;
        RECT 13.255 0.085 13.425 0.900 ;
        RECT 14.095 0.085 14.355 1.280 ;
        RECT 0.000 -0.085 14.720 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 10.725 2.635 10.895 2.805 ;
        RECT 11.185 2.635 11.355 2.805 ;
        RECT 11.645 2.635 11.815 2.805 ;
        RECT 12.105 2.635 12.275 2.805 ;
        RECT 12.565 2.635 12.735 2.805 ;
        RECT 13.025 2.635 13.195 2.805 ;
        RECT 13.485 2.635 13.655 2.805 ;
        RECT 13.945 2.635 14.115 2.805 ;
        RECT 14.405 2.635 14.575 2.805 ;
        RECT 0.635 1.785 0.805 1.955 ;
        RECT 1.015 1.445 1.185 1.615 ;
        RECT 1.355 0.425 1.525 0.595 ;
        RECT 3.805 0.765 3.975 0.935 ;
        RECT 7.510 1.785 7.680 1.955 ;
        RECT 4.185 0.425 4.355 0.595 ;
        RECT 4.615 0.425 4.785 0.595 ;
        RECT 7.100 1.445 7.270 1.615 ;
        RECT 6.530 0.425 6.700 0.595 ;
        RECT 10.100 1.785 10.270 1.955 ;
        RECT 10.520 1.445 10.690 1.615 ;
        RECT 12.000 0.765 12.170 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
        RECT 10.725 -0.085 10.895 0.085 ;
        RECT 11.185 -0.085 11.355 0.085 ;
        RECT 11.645 -0.085 11.815 0.085 ;
        RECT 12.105 -0.085 12.275 0.085 ;
        RECT 12.565 -0.085 12.735 0.085 ;
        RECT 13.025 -0.085 13.195 0.085 ;
        RECT 13.485 -0.085 13.655 0.085 ;
        RECT 13.945 -0.085 14.115 0.085 ;
        RECT 14.405 -0.085 14.575 0.085 ;
      LAYER met1 ;
        RECT 0.575 1.940 0.865 1.985 ;
        RECT 7.450 1.940 7.740 1.985 ;
        RECT 10.040 1.940 10.330 1.985 ;
        RECT 0.575 1.800 10.330 1.940 ;
        RECT 0.575 1.755 0.865 1.800 ;
        RECT 7.450 1.755 7.740 1.800 ;
        RECT 10.040 1.755 10.330 1.800 ;
        RECT 0.955 1.600 1.245 1.645 ;
        RECT 7.040 1.600 7.330 1.645 ;
        RECT 10.460 1.600 10.750 1.645 ;
        RECT 0.955 1.460 10.750 1.600 ;
        RECT 0.955 1.415 1.245 1.460 ;
        RECT 7.040 1.415 7.330 1.460 ;
        RECT 10.460 1.415 10.750 1.460 ;
        RECT 3.745 0.920 4.035 0.965 ;
        RECT 11.940 0.920 12.230 0.965 ;
        RECT 3.745 0.780 12.230 0.920 ;
        RECT 3.745 0.735 4.035 0.780 ;
        RECT 11.940 0.735 12.230 0.780 ;
        RECT 1.295 0.580 1.585 0.625 ;
        RECT 4.125 0.580 4.415 0.625 ;
        RECT 1.295 0.395 4.415 0.580 ;
        RECT 4.555 0.580 4.845 0.625 ;
        RECT 6.470 0.580 6.760 0.625 ;
        RECT 4.555 0.395 6.760 0.580 ;
  END
END sky130_fd_sc_hd__sedfxtp_4

#--------EOF---------

MACRO sky130_fd_sc_hd__tap_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tap_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.190 0.445 0.975 ;
      LAYER li1 ;
        RECT 0.085 0.265 0.375 0.810 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 2.910 ;
      LAYER li1 ;
        RECT 0.085 1.470 0.375 2.455 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.460 2.805 ;
        RECT 0.000 -0.085 0.460 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
  END
END sky130_fd_sc_hd__tap_1

#--------EOF---------

MACRO sky130_fd_sc_hd__tap_2
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tap_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.920 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 0.920 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.190 0.905 0.975 ;
      LAYER li1 ;
        RECT 0.085 0.265 0.835 0.810 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 1.110 2.910 ;
      LAYER li1 ;
        RECT 0.085 1.470 0.835 2.455 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.920 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.920 2.805 ;
        RECT 0.000 -0.085 0.920 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
  END
END sky130_fd_sc_hd__tap_2

#--------EOF---------

MACRO sky130_fd_sc_hd__tapvgnd2_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tapvgnd2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.190 0.445 0.975 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 2.910 ;
      LAYER met1 ;
        RECT 0.085 1.755 0.375 1.985 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.460 2.805 ;
        RECT 0.085 1.470 0.375 2.455 ;
        RECT 0.085 0.085 0.375 0.810 ;
        RECT 0.000 -0.085 0.460 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.145 1.785 0.315 1.955 ;
        RECT 0.145 -0.085 0.315 0.085 ;
  END
END sky130_fd_sc_hd__tapvgnd2_1

#--------EOF---------

MACRO sky130_fd_sc_hd__tapvgnd_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tapvgnd_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.190 0.445 0.975 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 2.910 ;
      LAYER met1 ;
        RECT 0.085 2.095 0.375 2.325 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.460 2.805 ;
        RECT 0.085 1.470 0.375 2.455 ;
        RECT 0.085 0.085 0.375 0.810 ;
        RECT 0.000 -0.085 0.460 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.145 2.125 0.315 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
  END
END sky130_fd_sc_hd__tapvgnd_1

#--------EOF---------

MACRO sky130_fd_sc_hd__tapvpwrvgnd_1
  CLASS CORE WELLTAP ;
  FOREIGN sky130_fd_sc_hd__tapvpwrvgnd_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.460 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER pwell ;
        RECT 0.015 0.190 0.445 0.975 ;
      LAYER met1 ;
        RECT 0.000 -0.240 0.460 0.240 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 0.650 2.910 ;
      LAYER met1 ;
        RECT 0.000 2.480 0.460 2.960 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 0.460 2.805 ;
        RECT 0.085 1.470 0.375 2.635 ;
        RECT 0.085 0.085 0.375 0.810 ;
        RECT 0.000 -0.085 0.460 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
  END
END sky130_fd_sc_hd__tapvpwrvgnd_1

#--------EOF---------

MACRO sky130_fd_sc_hd__xnor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.930 1.075 1.625 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.445 1.965 1.615 ;
        RECT 0.425 0.995 0.670 1.445 ;
        RECT 1.795 1.245 1.965 1.445 ;
        RECT 1.795 1.075 2.395 1.245 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.105 0.105 3.215 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.525000 ;
    PORT
      LAYER li1 ;
        RECT 2.265 2.125 2.645 2.295 ;
        RECT 2.475 1.955 2.645 2.125 ;
        RECT 2.475 1.755 3.135 1.955 ;
        RECT 2.965 0.825 3.135 1.755 ;
        RECT 2.815 0.345 3.135 0.825 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 2.125 0.385 2.635 ;
        RECT 0.555 1.955 0.885 2.465 ;
        RECT 1.055 2.125 1.685 2.635 ;
        RECT 2.815 2.125 3.115 2.635 ;
        RECT 0.085 1.785 2.305 1.955 ;
        RECT 0.085 0.825 0.255 1.785 ;
        RECT 2.135 1.585 2.305 1.785 ;
        RECT 2.135 1.415 2.795 1.585 ;
        RECT 2.625 0.995 2.795 1.415 ;
        RECT 0.085 0.280 0.550 0.825 ;
        RECT 1.055 0.085 1.225 0.905 ;
        RECT 1.395 0.825 2.305 0.905 ;
        RECT 1.395 0.735 2.645 0.825 ;
        RECT 1.395 0.255 1.725 0.735 ;
        RECT 2.135 0.655 2.645 0.735 ;
        RECT 1.895 0.085 2.245 0.475 ;
        RECT 2.415 0.255 2.645 0.655 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__xnor2_1

#--------EOF---------

MACRO sky130_fd_sc_hd__xnor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 1.255 1.075 2.705 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.790 1.445 3.100 1.615 ;
        RECT 0.790 1.285 0.960 1.445 ;
        RECT 0.485 1.075 0.960 1.285 ;
        RECT 2.930 1.285 3.100 1.445 ;
        RECT 2.930 1.075 3.955 1.285 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.845 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.913000 ;
    PORT
      LAYER li1 ;
        RECT 3.725 1.965 3.935 2.125 ;
        RECT 5.045 1.965 5.295 2.125 ;
        RECT 3.725 1.795 5.295 1.965 ;
        RECT 5.045 1.625 5.295 1.795 ;
        RECT 5.045 1.415 5.895 1.625 ;
        RECT 5.505 0.475 5.895 1.415 ;
        RECT 4.585 0.305 5.895 0.475 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.085 1.965 0.400 2.465 ;
        RECT 0.570 2.135 0.820 2.635 ;
        RECT 0.990 1.965 1.240 2.465 ;
        RECT 1.410 2.135 1.660 2.635 ;
        RECT 1.830 1.965 2.080 2.465 ;
        RECT 2.390 2.125 2.640 2.465 ;
        RECT 2.810 2.135 3.060 2.635 ;
        RECT 3.230 2.295 4.355 2.465 ;
        RECT 3.230 2.125 3.555 2.295 ;
        RECT 4.105 2.135 4.355 2.295 ;
        RECT 4.625 2.135 4.875 2.635 ;
        RECT 0.085 1.955 2.080 1.965 ;
        RECT 0.085 1.785 3.480 1.955 ;
        RECT 5.465 1.795 5.895 2.635 ;
        RECT 0.085 0.895 0.315 1.785 ;
        RECT 3.310 1.625 3.480 1.785 ;
        RECT 3.310 1.455 4.805 1.625 ;
        RECT 4.635 1.245 4.805 1.455 ;
        RECT 4.635 1.075 5.295 1.245 ;
        RECT 0.085 0.645 0.860 0.895 ;
        RECT 1.030 0.725 2.120 0.905 ;
        RECT 1.030 0.475 1.280 0.725 ;
        RECT 0.105 0.255 1.280 0.475 ;
        RECT 1.450 0.085 1.620 0.555 ;
        RECT 1.790 0.255 2.120 0.725 ;
        RECT 2.430 0.085 2.600 0.905 ;
        RECT 2.770 0.725 5.335 0.905 ;
        RECT 2.770 0.255 3.100 0.725 ;
        RECT 3.270 0.085 3.440 0.555 ;
        RECT 3.610 0.255 3.975 0.725 ;
        RECT 5.005 0.645 5.335 0.725 ;
        RECT 4.145 0.085 4.315 0.555 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 2.465 2.125 2.635 2.295 ;
        RECT 3.385 2.125 3.555 2.295 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
      LAYER met1 ;
        RECT 2.405 2.280 2.695 2.325 ;
        RECT 3.325 2.280 3.615 2.325 ;
        RECT 2.405 2.140 3.615 2.280 ;
        RECT 2.405 2.095 2.695 2.140 ;
        RECT 3.325 2.095 3.615 2.140 ;
  END
END sky130_fd_sc_hd__xnor2_2

#--------EOF---------

MACRO sky130_fd_sc_hd__xnor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 2.175 1.075 5.390 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 1.685 1.445 5.730 1.615 ;
        RECT 1.685 1.275 1.855 1.445 ;
        RECT 0.490 1.075 1.855 1.275 ;
        RECT 5.560 1.275 5.730 1.445 ;
        RECT 5.560 1.075 7.430 1.275 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.060 0.105 10.080 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.721000 ;
    PORT
      LAYER li1 ;
        RECT 7.960 2.045 8.250 2.465 ;
        RECT 6.160 1.785 8.250 2.045 ;
        RECT 7.960 1.665 8.250 1.785 ;
        RECT 8.840 1.665 9.090 2.465 ;
        RECT 9.680 1.665 10.035 2.465 ;
        RECT 7.960 1.445 10.035 1.665 ;
        RECT 9.815 0.905 10.035 1.445 ;
        RECT 8.380 0.645 10.035 0.905 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.085 1.615 0.460 2.465 ;
        RECT 0.630 1.835 0.880 2.635 ;
        RECT 1.050 2.005 1.300 2.465 ;
        RECT 1.470 2.175 1.720 2.635 ;
        RECT 1.890 2.005 2.140 2.465 ;
        RECT 2.310 2.175 2.560 2.635 ;
        RECT 2.730 2.005 2.980 2.465 ;
        RECT 3.150 2.175 3.400 2.635 ;
        RECT 3.570 2.005 3.820 2.465 ;
        RECT 1.050 1.785 3.820 2.005 ;
        RECT 4.035 2.005 4.350 2.465 ;
        RECT 4.520 2.175 4.770 2.635 ;
        RECT 4.940 2.005 5.190 2.465 ;
        RECT 5.360 2.175 5.610 2.635 ;
        RECT 5.780 2.215 7.750 2.465 ;
        RECT 5.780 2.005 5.990 2.215 ;
        RECT 4.035 1.785 5.990 2.005 ;
        RECT 8.420 1.835 8.670 2.635 ;
        RECT 9.260 1.835 9.510 2.635 ;
        RECT 1.050 1.615 1.300 1.785 ;
        RECT 0.085 1.445 1.300 1.615 ;
        RECT 5.900 1.445 7.770 1.615 ;
        RECT 0.085 0.905 0.320 1.445 ;
        RECT 7.600 1.275 7.770 1.445 ;
        RECT 7.600 1.075 9.645 1.275 ;
        RECT 0.085 0.645 1.760 0.905 ;
        RECT 1.930 0.725 3.860 0.905 ;
        RECT 1.930 0.475 2.180 0.725 ;
        RECT 0.170 0.255 2.180 0.475 ;
        RECT 2.350 0.085 2.520 0.555 ;
        RECT 2.690 0.255 3.020 0.725 ;
        RECT 3.190 0.085 3.360 0.555 ;
        RECT 3.530 0.255 3.860 0.725 ;
        RECT 4.035 0.085 4.310 0.905 ;
        RECT 4.480 0.735 8.210 0.905 ;
        RECT 4.480 0.725 7.430 0.735 ;
        RECT 4.480 0.255 4.810 0.725 ;
        RECT 4.980 0.085 5.150 0.555 ;
        RECT 5.320 0.255 5.650 0.725 ;
        RECT 5.820 0.085 5.990 0.555 ;
        RECT 6.160 0.255 6.490 0.725 ;
        RECT 6.660 0.085 6.830 0.555 ;
        RECT 7.000 0.255 7.330 0.725 ;
        RECT 7.500 0.085 7.770 0.555 ;
        RECT 7.960 0.475 8.210 0.735 ;
        RECT 7.960 0.305 9.970 0.475 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 1.065 1.445 1.235 1.615 ;
        RECT 6.125 1.445 6.295 1.615 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
      LAYER met1 ;
        RECT 1.005 1.600 1.295 1.645 ;
        RECT 6.065 1.600 6.355 1.645 ;
        RECT 1.005 1.460 6.355 1.600 ;
        RECT 1.005 1.415 1.295 1.460 ;
        RECT 6.065 1.415 6.355 1.460 ;
  END
END sky130_fd_sc_hd__xnor2_4

#--------EOF---------

MACRO sky130_fd_sc_hd__xnor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 7.045 1.075 7.455 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.661500 ;
    PORT
      LAYER li1 ;
        RECT 6.225 1.445 6.805 1.615 ;
        RECT 6.225 0.995 6.395 1.445 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.381000 ;
    PORT
      LAYER li1 ;
        RECT 1.615 1.075 2.180 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.005 6.705 1.015 ;
        RECT 0.005 0.115 8.260 1.005 ;
        RECT 0.005 0.105 0.985 0.115 ;
        RECT 3.275 0.105 4.225 0.115 ;
        RECT 6.280 0.105 8.260 0.115 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.470 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.449000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.440 0.365 2.465 ;
        RECT 0.085 0.925 0.330 1.440 ;
        RECT 0.085 0.350 0.345 0.925 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.280 2.805 ;
        RECT 0.535 2.215 0.870 2.635 ;
        RECT 1.050 2.235 2.520 2.405 ;
        RECT 3.225 2.235 3.555 2.635 ;
        RECT 3.890 2.275 6.985 2.445 ;
        RECT 7.395 2.275 7.730 2.635 ;
        RECT 1.050 2.045 1.220 2.235 ;
        RECT 3.890 2.065 4.060 2.275 ;
        RECT 0.535 1.875 1.220 2.045 ;
        RECT 1.560 1.895 4.060 2.065 ;
        RECT 0.535 1.325 0.705 1.875 ;
        RECT 0.935 1.535 2.520 1.705 ;
        RECT 0.500 0.995 0.705 1.325 ;
        RECT 0.530 0.865 0.705 0.995 ;
        RECT 0.530 0.695 1.105 0.865 ;
        RECT 0.515 0.085 0.765 0.525 ;
        RECT 0.935 0.425 1.105 0.695 ;
        RECT 1.275 0.595 1.445 1.535 ;
        RECT 2.350 1.325 2.520 1.535 ;
        RECT 2.690 1.525 3.075 1.695 ;
        RECT 2.795 1.375 3.075 1.525 ;
        RECT 2.350 0.995 2.625 1.325 ;
        RECT 1.745 0.795 2.125 0.905 ;
        RECT 2.795 0.795 2.965 1.375 ;
        RECT 3.245 1.205 3.415 1.895 ;
        RECT 3.645 1.445 4.065 1.715 ;
        RECT 1.745 0.625 2.965 0.795 ;
        RECT 3.135 1.035 3.415 1.205 ;
        RECT 3.135 0.455 3.305 1.035 ;
        RECT 2.070 0.425 2.505 0.455 ;
        RECT 0.935 0.255 2.505 0.425 ;
        RECT 2.675 0.285 3.305 0.455 ;
        RECT 3.475 0.085 3.645 0.865 ;
        RECT 3.825 0.415 4.065 1.445 ;
        RECT 4.245 0.595 4.415 2.105 ;
        RECT 4.585 0.890 4.755 2.275 ;
        RECT 7.900 2.105 8.195 2.465 ;
        RECT 4.935 1.615 5.350 2.045 ;
        RECT 5.885 1.935 8.195 2.105 ;
        RECT 4.935 1.445 5.715 1.615 ;
        RECT 4.950 0.995 5.375 1.270 ;
        RECT 4.585 0.825 4.795 0.890 ;
        RECT 4.585 0.720 4.995 0.825 ;
        RECT 4.625 0.655 4.995 0.720 ;
        RECT 4.245 0.485 4.455 0.595 ;
        RECT 4.245 0.265 4.655 0.485 ;
        RECT 4.825 0.320 4.995 0.655 ;
        RECT 5.165 0.630 5.375 0.995 ;
        RECT 5.545 0.425 5.715 1.445 ;
        RECT 5.885 0.595 6.055 1.935 ;
        RECT 7.710 1.875 8.195 1.935 ;
        RECT 6.975 1.495 7.795 1.705 ;
        RECT 7.625 1.325 7.795 1.495 ;
        RECT 6.565 0.945 6.875 1.275 ;
        RECT 7.625 0.995 7.855 1.325 ;
        RECT 6.565 0.730 6.770 0.945 ;
        RECT 7.625 0.905 7.795 0.995 ;
        RECT 7.055 0.750 7.795 0.905 ;
        RECT 7.015 0.735 7.795 0.750 ;
        RECT 6.225 0.425 6.690 0.465 ;
        RECT 5.545 0.255 6.690 0.425 ;
        RECT 7.015 0.295 7.305 0.735 ;
        RECT 8.025 0.585 8.195 1.875 ;
        RECT 7.475 0.085 7.645 0.565 ;
        RECT 7.895 0.255 8.195 0.585 ;
        RECT 0.000 -0.085 8.280 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 2.905 1.445 3.075 1.615 ;
        RECT 3.825 0.765 3.995 0.935 ;
        RECT 5.205 1.445 5.375 1.615 ;
        RECT 4.285 0.425 4.455 0.595 ;
        RECT 5.205 0.765 5.375 0.935 ;
        RECT 6.585 0.765 6.755 0.935 ;
        RECT 7.045 0.425 7.215 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
      LAYER met1 ;
        RECT 2.845 1.600 3.135 1.645 ;
        RECT 5.145 1.600 5.435 1.645 ;
        RECT 2.845 1.460 5.435 1.600 ;
        RECT 2.845 1.415 3.135 1.460 ;
        RECT 5.145 1.415 5.435 1.460 ;
        RECT 3.765 0.920 4.055 0.965 ;
        RECT 5.145 0.920 5.435 0.965 ;
        RECT 6.525 0.920 6.815 0.965 ;
        RECT 3.765 0.780 6.815 0.920 ;
        RECT 3.765 0.735 4.055 0.780 ;
        RECT 5.145 0.735 5.435 0.780 ;
        RECT 6.525 0.735 6.815 0.780 ;
        RECT 4.225 0.580 4.515 0.625 ;
        RECT 6.985 0.580 7.275 0.625 ;
        RECT 4.225 0.440 7.275 0.580 ;
        RECT 4.225 0.395 4.515 0.440 ;
        RECT 6.985 0.395 7.275 0.440 ;
  END
END sky130_fd_sc_hd__xnor3_1

#--------EOF---------

MACRO sky130_fd_sc_hd__xnor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 7.505 1.075 7.915 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.661500 ;
    PORT
      LAYER li1 ;
        RECT 6.685 1.445 7.265 1.615 ;
        RECT 6.685 0.995 6.855 1.445 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.381000 ;
    PORT
      LAYER li1 ;
        RECT 2.075 1.075 2.640 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.005 7.165 1.015 ;
        RECT 0.005 0.115 8.720 1.005 ;
        RECT 0.005 0.105 1.445 0.115 ;
        RECT 3.735 0.105 4.685 0.115 ;
        RECT 6.740 0.105 8.720 0.115 ;
        RECT 0.150 -0.085 0.320 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.545 1.440 0.825 2.465 ;
        RECT 0.545 0.925 0.790 1.440 ;
        RECT 0.545 0.350 0.805 0.925 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.740 2.805 ;
        RECT 0.085 1.490 0.375 2.635 ;
        RECT 0.995 2.215 1.330 2.635 ;
        RECT 1.510 2.235 2.980 2.405 ;
        RECT 3.685 2.235 4.015 2.635 ;
        RECT 4.350 2.275 7.445 2.445 ;
        RECT 7.855 2.275 8.190 2.635 ;
        RECT 1.510 2.045 1.680 2.235 ;
        RECT 4.350 2.065 4.520 2.275 ;
        RECT 0.995 1.875 1.680 2.045 ;
        RECT 2.020 1.895 4.520 2.065 ;
        RECT 0.995 1.325 1.165 1.875 ;
        RECT 1.395 1.535 2.980 1.705 ;
        RECT 0.960 0.995 1.165 1.325 ;
        RECT 0.990 0.865 1.165 0.995 ;
        RECT 0.085 0.085 0.375 0.735 ;
        RECT 0.990 0.695 1.565 0.865 ;
        RECT 0.975 0.085 1.225 0.525 ;
        RECT 1.395 0.425 1.565 0.695 ;
        RECT 1.735 0.595 1.905 1.535 ;
        RECT 2.810 1.325 2.980 1.535 ;
        RECT 3.150 1.525 3.535 1.695 ;
        RECT 3.255 1.375 3.535 1.525 ;
        RECT 2.810 0.995 3.085 1.325 ;
        RECT 2.205 0.795 2.585 0.905 ;
        RECT 3.255 0.795 3.425 1.375 ;
        RECT 3.705 1.205 3.875 1.895 ;
        RECT 4.105 1.445 4.525 1.715 ;
        RECT 2.205 0.625 3.425 0.795 ;
        RECT 3.595 1.035 3.875 1.205 ;
        RECT 3.595 0.455 3.765 1.035 ;
        RECT 2.530 0.425 2.965 0.455 ;
        RECT 1.395 0.255 2.965 0.425 ;
        RECT 3.135 0.285 3.765 0.455 ;
        RECT 3.935 0.085 4.105 0.865 ;
        RECT 4.285 0.415 4.525 1.445 ;
        RECT 4.705 0.595 4.875 2.105 ;
        RECT 5.045 0.890 5.215 2.275 ;
        RECT 8.360 2.105 8.655 2.465 ;
        RECT 5.395 1.615 5.810 2.045 ;
        RECT 6.345 1.935 8.655 2.105 ;
        RECT 5.395 1.445 6.175 1.615 ;
        RECT 5.410 0.995 5.835 1.270 ;
        RECT 5.045 0.825 5.255 0.890 ;
        RECT 5.045 0.720 5.455 0.825 ;
        RECT 5.085 0.655 5.455 0.720 ;
        RECT 4.705 0.485 4.915 0.595 ;
        RECT 4.705 0.265 5.115 0.485 ;
        RECT 5.285 0.320 5.455 0.655 ;
        RECT 5.625 0.630 5.835 0.995 ;
        RECT 6.005 0.425 6.175 1.445 ;
        RECT 6.345 0.595 6.515 1.935 ;
        RECT 8.170 1.875 8.655 1.935 ;
        RECT 7.435 1.495 8.255 1.705 ;
        RECT 8.085 1.325 8.255 1.495 ;
        RECT 7.025 0.945 7.335 1.275 ;
        RECT 8.085 0.995 8.315 1.325 ;
        RECT 7.025 0.730 7.230 0.945 ;
        RECT 8.085 0.905 8.255 0.995 ;
        RECT 7.515 0.750 8.255 0.905 ;
        RECT 7.475 0.735 8.255 0.750 ;
        RECT 6.685 0.425 7.150 0.465 ;
        RECT 6.005 0.255 7.150 0.425 ;
        RECT 7.475 0.295 7.765 0.735 ;
        RECT 8.485 0.585 8.655 1.875 ;
        RECT 7.935 0.085 8.105 0.565 ;
        RECT 8.355 0.255 8.655 0.585 ;
        RECT 0.000 -0.085 8.740 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 3.365 1.445 3.535 1.615 ;
        RECT 4.285 0.765 4.455 0.935 ;
        RECT 5.665 1.445 5.835 1.615 ;
        RECT 4.745 0.425 4.915 0.595 ;
        RECT 5.665 0.765 5.835 0.935 ;
        RECT 7.045 0.765 7.215 0.935 ;
        RECT 7.505 0.425 7.675 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
      LAYER met1 ;
        RECT 3.305 1.600 3.595 1.645 ;
        RECT 5.605 1.600 5.895 1.645 ;
        RECT 3.305 1.460 5.895 1.600 ;
        RECT 3.305 1.415 3.595 1.460 ;
        RECT 5.605 1.415 5.895 1.460 ;
        RECT 4.225 0.920 4.515 0.965 ;
        RECT 5.605 0.920 5.895 0.965 ;
        RECT 6.985 0.920 7.275 0.965 ;
        RECT 4.225 0.780 7.275 0.920 ;
        RECT 4.225 0.735 4.515 0.780 ;
        RECT 5.605 0.735 5.895 0.780 ;
        RECT 6.985 0.735 7.275 0.780 ;
        RECT 4.685 0.580 4.975 0.625 ;
        RECT 7.445 0.580 7.735 0.625 ;
        RECT 4.685 0.440 7.735 0.580 ;
        RECT 4.685 0.395 4.975 0.440 ;
        RECT 7.445 0.395 7.735 0.440 ;
  END
END sky130_fd_sc_hd__xnor3_2

#--------EOF---------

MACRO sky130_fd_sc_hd__xnor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xnor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 8.425 1.075 8.835 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.661500 ;
    PORT
      LAYER li1 ;
        RECT 7.605 1.445 8.185 1.615 ;
        RECT 7.605 0.995 7.775 1.445 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.381000 ;
    PORT
      LAYER li1 ;
        RECT 2.995 1.075 3.560 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.115 1.005 8.085 1.015 ;
        RECT 0.115 0.115 9.640 1.005 ;
        RECT 0.115 0.105 2.365 0.115 ;
        RECT 4.655 0.105 5.605 0.115 ;
        RECT 7.660 0.105 9.640 0.115 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.625 1.325 0.955 2.425 ;
        RECT 1.465 1.440 1.745 2.465 ;
        RECT 1.465 1.325 1.710 1.440 ;
        RECT 0.625 0.995 1.710 1.325 ;
        RECT 0.625 0.375 0.875 0.995 ;
        RECT 1.465 0.925 1.710 0.995 ;
        RECT 1.465 0.350 1.725 0.925 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 0.285 1.490 0.455 2.635 ;
        RECT 1.125 1.495 1.295 2.635 ;
        RECT 1.915 2.215 2.250 2.635 ;
        RECT 2.430 2.235 3.900 2.405 ;
        RECT 4.605 2.235 4.935 2.635 ;
        RECT 5.270 2.275 8.365 2.445 ;
        RECT 8.775 2.275 9.110 2.635 ;
        RECT 2.430 2.045 2.600 2.235 ;
        RECT 5.270 2.065 5.440 2.275 ;
        RECT 1.915 1.875 2.600 2.045 ;
        RECT 2.940 1.895 5.440 2.065 ;
        RECT 1.915 1.325 2.085 1.875 ;
        RECT 2.315 1.535 3.900 1.705 ;
        RECT 1.880 0.995 2.085 1.325 ;
        RECT 1.910 0.865 2.085 0.995 ;
        RECT 0.285 0.085 0.455 0.735 ;
        RECT 1.125 0.085 1.295 0.735 ;
        RECT 1.910 0.695 2.485 0.865 ;
        RECT 1.895 0.085 2.145 0.525 ;
        RECT 2.315 0.425 2.485 0.695 ;
        RECT 2.655 0.595 2.825 1.535 ;
        RECT 3.730 1.325 3.900 1.535 ;
        RECT 4.070 1.525 4.455 1.695 ;
        RECT 4.175 1.375 4.455 1.525 ;
        RECT 3.730 0.995 4.005 1.325 ;
        RECT 3.125 0.795 3.505 0.905 ;
        RECT 4.175 0.795 4.345 1.375 ;
        RECT 4.625 1.205 4.795 1.895 ;
        RECT 5.025 1.445 5.445 1.715 ;
        RECT 3.125 0.625 4.345 0.795 ;
        RECT 4.515 1.035 4.795 1.205 ;
        RECT 4.515 0.455 4.685 1.035 ;
        RECT 3.450 0.425 3.885 0.455 ;
        RECT 2.315 0.255 3.885 0.425 ;
        RECT 4.055 0.285 4.685 0.455 ;
        RECT 4.855 0.085 5.025 0.865 ;
        RECT 5.205 0.415 5.445 1.445 ;
        RECT 5.625 0.595 5.795 2.105 ;
        RECT 5.965 0.890 6.135 2.275 ;
        RECT 9.280 2.105 9.575 2.465 ;
        RECT 6.315 1.615 6.730 2.045 ;
        RECT 7.265 1.935 9.575 2.105 ;
        RECT 6.315 1.445 7.095 1.615 ;
        RECT 6.330 0.995 6.755 1.270 ;
        RECT 5.965 0.825 6.175 0.890 ;
        RECT 5.965 0.720 6.375 0.825 ;
        RECT 6.005 0.655 6.375 0.720 ;
        RECT 5.625 0.485 5.835 0.595 ;
        RECT 5.625 0.265 6.035 0.485 ;
        RECT 6.205 0.320 6.375 0.655 ;
        RECT 6.545 0.630 6.755 0.995 ;
        RECT 6.925 0.425 7.095 1.445 ;
        RECT 7.265 0.595 7.435 1.935 ;
        RECT 9.090 1.875 9.575 1.935 ;
        RECT 8.355 1.495 9.175 1.705 ;
        RECT 9.005 1.325 9.175 1.495 ;
        RECT 7.945 0.945 8.255 1.275 ;
        RECT 9.005 0.995 9.235 1.325 ;
        RECT 7.945 0.730 8.150 0.945 ;
        RECT 9.005 0.905 9.175 0.995 ;
        RECT 8.435 0.750 9.175 0.905 ;
        RECT 8.395 0.735 9.175 0.750 ;
        RECT 7.605 0.425 8.070 0.465 ;
        RECT 6.925 0.255 8.070 0.425 ;
        RECT 8.395 0.295 8.685 0.735 ;
        RECT 9.405 0.585 9.575 1.875 ;
        RECT 8.855 0.085 9.025 0.565 ;
        RECT 9.275 0.255 9.575 0.585 ;
        RECT 0.000 -0.085 9.660 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 4.285 1.445 4.455 1.615 ;
        RECT 5.205 0.765 5.375 0.935 ;
        RECT 6.585 1.445 6.755 1.615 ;
        RECT 5.665 0.425 5.835 0.595 ;
        RECT 6.585 0.765 6.755 0.935 ;
        RECT 7.965 0.765 8.135 0.935 ;
        RECT 8.425 0.425 8.595 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 4.225 1.600 4.515 1.645 ;
        RECT 6.525 1.600 6.815 1.645 ;
        RECT 4.225 1.460 6.815 1.600 ;
        RECT 4.225 1.415 4.515 1.460 ;
        RECT 6.525 1.415 6.815 1.460 ;
        RECT 5.145 0.920 5.435 0.965 ;
        RECT 6.525 0.920 6.815 0.965 ;
        RECT 7.905 0.920 8.195 0.965 ;
        RECT 5.145 0.780 8.195 0.920 ;
        RECT 5.145 0.735 5.435 0.780 ;
        RECT 6.525 0.735 6.815 0.780 ;
        RECT 7.905 0.735 8.195 0.780 ;
        RECT 5.605 0.580 5.895 0.625 ;
        RECT 8.365 0.580 8.655 0.625 ;
        RECT 5.605 0.440 8.655 0.580 ;
        RECT 5.605 0.395 5.895 0.440 ;
        RECT 8.365 0.395 8.655 0.440 ;
  END
END sky130_fd_sc_hd__xnor3_4

#--------EOF---------

MACRO sky130_fd_sc_hd__xor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor2_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.220 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.840 1.075 1.390 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER li1 ;
        RECT 0.425 1.445 1.730 1.615 ;
        RECT 0.425 0.995 0.670 1.445 ;
        RECT 1.560 1.245 1.730 1.445 ;
        RECT 1.560 1.075 1.935 1.245 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 3.220 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.045 0.105 3.215 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 3.410 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 3.220 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.800500 ;
    PORT
      LAYER li1 ;
        RECT 2.815 1.535 3.135 2.465 ;
        RECT 2.505 1.365 3.135 1.535 ;
        RECT 2.505 0.485 2.675 1.365 ;
        RECT 1.720 0.315 2.675 0.485 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 3.220 2.805 ;
        RECT 0.085 1.785 0.465 2.465 ;
        RECT 1.055 1.785 1.225 2.635 ;
        RECT 1.395 1.955 1.725 2.465 ;
        RECT 1.895 2.125 2.065 2.635 ;
        RECT 2.235 1.955 2.635 2.465 ;
        RECT 1.395 1.785 2.635 1.955 ;
        RECT 0.085 0.825 0.255 1.785 ;
        RECT 2.105 0.825 2.335 1.325 ;
        RECT 0.085 0.655 2.335 0.825 ;
        RECT 0.135 0.085 0.465 0.475 ;
        RECT 0.635 0.335 0.805 0.655 ;
        RECT 0.975 0.085 1.305 0.475 ;
        RECT 2.845 0.085 3.135 0.920 ;
        RECT 0.000 -0.085 3.220 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
  END
END sky130_fd_sc_hd__xor2_1

#--------EOF---------

MACRO sky130_fd_sc_hd__xor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor2_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.980 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER li1 ;
        RECT 0.705 1.445 1.880 1.615 ;
        RECT 0.705 1.275 0.875 1.445 ;
        RECT 0.545 1.075 0.875 1.275 ;
        RECT 1.710 1.275 1.880 1.445 ;
        RECT 1.710 1.075 3.230 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met1 ;
        RECT 1.005 1.260 1.295 1.305 ;
        RECT 3.765 1.260 4.055 1.305 ;
        RECT 1.005 1.120 4.055 1.260 ;
        RECT 1.005 1.075 1.295 1.120 ;
        RECT 3.765 1.075 4.055 1.120 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.980 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.825 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 6.170 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.980 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.656750 ;
    PORT
      LAYER li1 ;
        RECT 5.025 1.625 5.275 2.125 ;
        RECT 5.025 1.415 5.895 1.625 ;
        RECT 5.485 0.905 5.895 1.415 ;
        RECT 3.625 0.725 5.895 0.905 ;
        RECT 3.625 0.645 3.955 0.725 ;
        RECT 4.985 0.645 5.315 0.725 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 5.980 2.805 ;
        RECT 0.120 2.135 0.400 2.465 ;
        RECT 0.570 2.135 0.820 2.635 ;
        RECT 0.990 2.295 2.080 2.465 ;
        RECT 0.990 2.135 1.240 2.295 ;
        RECT 1.830 2.135 2.080 2.295 ;
        RECT 0.145 2.125 0.315 2.135 ;
        RECT 1.065 2.125 1.235 2.135 ;
        RECT 2.285 2.125 2.600 2.465 ;
        RECT 2.770 2.135 3.020 2.635 ;
        RECT 1.410 1.955 1.660 2.125 ;
        RECT 2.390 1.955 2.600 2.125 ;
        RECT 3.190 1.955 3.440 2.465 ;
        RECT 3.610 2.135 3.915 2.635 ;
        RECT 4.085 2.295 5.695 2.465 ;
        RECT 4.085 1.955 4.855 2.295 ;
        RECT 0.120 1.785 2.220 1.955 ;
        RECT 2.390 1.785 4.855 1.955 ;
        RECT 5.445 1.795 5.695 2.295 ;
        RECT 0.120 0.905 0.290 1.785 ;
        RECT 2.050 1.615 2.220 1.785 ;
        RECT 2.050 1.445 4.785 1.615 ;
        RECT 1.045 1.075 1.540 1.275 ;
        RECT 3.420 1.075 4.090 1.275 ;
        RECT 4.615 1.245 4.785 1.445 ;
        RECT 4.615 1.075 5.275 1.245 ;
        RECT 0.120 0.725 1.700 0.905 ;
        RECT 0.190 0.085 0.360 0.555 ;
        RECT 0.530 0.255 0.860 0.725 ;
        RECT 1.030 0.085 1.200 0.555 ;
        RECT 1.370 0.255 1.700 0.725 ;
        RECT 2.310 0.725 3.400 0.905 ;
        RECT 1.870 0.085 2.040 0.555 ;
        RECT 2.310 0.255 2.640 0.725 ;
        RECT 2.810 0.085 2.980 0.555 ;
        RECT 3.150 0.475 3.400 0.725 ;
        RECT 3.150 0.255 4.380 0.475 ;
        RECT 4.645 0.085 4.815 0.555 ;
        RECT 5.485 0.085 5.655 0.555 ;
        RECT 0.000 -0.085 5.980 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 1.065 1.105 1.235 1.275 ;
        RECT 3.825 1.105 3.995 1.275 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
      LAYER met1 ;
        RECT 0.085 2.280 0.375 2.325 ;
        RECT 1.005 2.280 1.295 2.325 ;
        RECT 0.085 2.140 1.295 2.280 ;
        RECT 0.085 2.095 0.375 2.140 ;
        RECT 1.005 2.095 1.295 2.140 ;
  END
END sky130_fd_sc_hd__xor2_2

#--------EOF---------

MACRO sky130_fd_sc_hd__xor2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor2_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 2.630 1.445 6.165 1.615 ;
        RECT 2.630 1.275 2.800 1.445 ;
        RECT 0.425 1.075 2.800 1.275 ;
        RECT 5.995 1.275 6.165 1.445 ;
        RECT 5.995 1.075 7.370 1.275 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.980000 ;
    PORT
      LAYER li1 ;
        RECT 2.970 1.105 5.740 1.275 ;
        RECT 2.970 1.075 5.000 1.105 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 10.000 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.524450 ;
    PORT
      LAYER met1 ;
        RECT 5.145 0.920 5.435 0.965 ;
        RECT 7.905 0.920 8.195 0.965 ;
        RECT 5.145 0.780 8.195 0.920 ;
        RECT 5.145 0.735 5.435 0.780 ;
        RECT 7.905 0.735 8.195 0.780 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.085 2.005 0.400 2.465 ;
        RECT 0.570 2.175 0.820 2.635 ;
        RECT 0.990 2.005 1.240 2.465 ;
        RECT 1.410 2.175 1.660 2.635 ;
        RECT 1.830 2.295 3.760 2.465 ;
        RECT 1.830 2.005 2.080 2.295 ;
        RECT 2.670 2.125 2.920 2.295 ;
        RECT 0.085 1.785 2.080 2.005 ;
        RECT 2.250 1.955 2.500 2.125 ;
        RECT 3.090 1.955 3.340 2.125 ;
        RECT 2.250 1.785 3.340 1.955 ;
        RECT 3.510 1.795 3.760 2.295 ;
        RECT 4.030 2.005 4.280 2.465 ;
        RECT 4.450 2.175 4.700 2.635 ;
        RECT 4.870 2.005 5.120 2.465 ;
        RECT 5.290 2.175 5.540 2.635 ;
        RECT 5.710 2.005 5.960 2.465 ;
        RECT 6.130 2.175 6.380 2.635 ;
        RECT 6.550 2.005 6.800 2.465 ;
        RECT 6.970 2.175 7.220 2.635 ;
        RECT 7.390 2.295 9.430 2.465 ;
        RECT 7.390 2.005 7.640 2.295 ;
        RECT 4.030 1.785 7.640 2.005 ;
        RECT 2.250 1.615 2.420 1.785 ;
        RECT 0.085 1.445 2.420 1.615 ;
        RECT 6.550 1.455 6.800 1.785 ;
        RECT 7.880 1.665 8.170 2.125 ;
        RECT 8.340 1.835 8.590 2.295 ;
        RECT 8.760 1.665 9.010 2.125 ;
        RECT 9.180 1.795 9.430 2.295 ;
        RECT 7.880 1.625 9.010 1.665 ;
        RECT 9.600 1.625 10.035 2.465 ;
        RECT 7.260 1.445 7.710 1.615 ;
        RECT 7.880 1.445 10.035 1.625 ;
        RECT 0.085 0.905 0.255 1.445 ;
        RECT 7.540 1.275 7.710 1.445 ;
        RECT 7.540 1.105 9.565 1.275 ;
        RECT 8.540 1.075 9.565 1.105 ;
        RECT 5.150 0.905 5.580 0.935 ;
        RECT 7.850 0.905 8.305 0.935 ;
        RECT 9.735 0.905 10.035 1.445 ;
        RECT 0.085 0.735 3.380 0.905 ;
        RECT 0.530 0.725 3.380 0.735 ;
        RECT 0.085 0.085 0.360 0.565 ;
        RECT 0.530 0.255 0.860 0.725 ;
        RECT 1.030 0.085 1.200 0.555 ;
        RECT 1.370 0.255 1.700 0.725 ;
        RECT 1.870 0.085 2.040 0.555 ;
        RECT 2.210 0.255 2.540 0.725 ;
        RECT 2.710 0.085 2.880 0.555 ;
        RECT 3.050 0.255 3.380 0.725 ;
        RECT 3.550 0.085 3.820 0.895 ;
        RECT 4.165 0.645 5.580 0.905 ;
        RECT 5.750 0.725 7.680 0.905 ;
        RECT 7.850 0.735 10.035 0.905 ;
        RECT 7.850 0.725 8.630 0.735 ;
        RECT 5.750 0.475 6.000 0.725 ;
        RECT 3.990 0.255 6.000 0.475 ;
        RECT 6.170 0.085 6.340 0.555 ;
        RECT 6.510 0.255 6.840 0.725 ;
        RECT 7.010 0.085 7.180 0.555 ;
        RECT 7.350 0.255 7.680 0.725 ;
        RECT 7.960 0.085 8.130 0.555 ;
        RECT 8.300 0.255 8.630 0.725 ;
        RECT 8.800 0.085 8.970 0.555 ;
        RECT 9.140 0.255 9.470 0.735 ;
        RECT 9.640 0.085 9.810 0.555 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 1.985 1.445 2.155 1.615 ;
        RECT 7.505 1.445 7.675 1.615 ;
        RECT 5.205 0.765 5.375 0.935 ;
        RECT 7.965 0.765 8.135 0.935 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
      LAYER met1 ;
        RECT 1.925 1.600 2.215 1.645 ;
        RECT 7.445 1.600 7.735 1.645 ;
        RECT 1.925 1.460 7.735 1.600 ;
        RECT 1.925 1.415 2.215 1.460 ;
        RECT 7.445 1.415 7.735 1.460 ;
  END
END sky130_fd_sc_hd__xor2_4

#--------EOF---------

MACRO sky130_fd_sc_hd__xor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor3_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.740 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 7.505 1.075 7.915 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.661500 ;
    PORT
      LAYER li1 ;
        RECT 6.685 1.445 7.265 1.615 ;
        RECT 6.685 0.995 6.855 1.445 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.381000 ;
    PORT
      LAYER li1 ;
        RECT 1.860 0.995 2.495 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.740 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.170 1.005 7.165 1.015 ;
        RECT 0.170 0.115 8.720 1.005 ;
        RECT 0.170 0.105 1.235 0.115 ;
        RECT 3.720 0.105 4.680 0.115 ;
        RECT 6.740 0.105 8.720 0.115 ;
        RECT 0.170 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 8.930 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.740 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.449000 ;
    PORT
      LAYER li1 ;
        RECT 0.085 1.440 0.610 2.465 ;
        RECT 0.085 0.925 0.400 1.440 ;
        RECT 0.085 0.350 0.590 0.925 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 8.740 2.805 ;
        RECT 0.780 2.215 1.115 2.635 ;
        RECT 1.300 2.235 2.895 2.405 ;
        RECT 3.110 2.235 3.515 2.405 ;
        RECT 3.685 2.235 4.015 2.635 ;
        RECT 4.350 2.275 7.445 2.445 ;
        RECT 7.855 2.275 8.190 2.635 ;
        RECT 1.300 2.045 1.470 2.235 ;
        RECT 3.345 2.065 3.515 2.235 ;
        RECT 4.350 2.065 4.520 2.275 ;
        RECT 0.780 1.875 1.470 2.045 ;
        RECT 1.870 1.895 3.175 2.065 ;
        RECT 3.345 1.895 4.520 2.065 ;
        RECT 0.780 1.325 0.950 1.875 ;
        RECT 1.185 1.535 2.835 1.705 ;
        RECT 0.750 0.995 0.950 1.325 ;
        RECT 0.780 0.865 0.950 0.995 ;
        RECT 0.780 0.695 1.350 0.865 ;
        RECT 0.760 0.085 1.010 0.525 ;
        RECT 1.180 0.425 1.350 0.695 ;
        RECT 1.520 0.595 1.690 1.535 ;
        RECT 2.665 1.325 2.835 1.535 ;
        RECT 3.005 1.695 3.175 1.895 ;
        RECT 3.005 1.525 3.535 1.695 ;
        RECT 3.250 1.375 3.535 1.525 ;
        RECT 2.665 0.995 2.940 1.325 ;
        RECT 1.970 0.655 3.080 0.825 ;
        RECT 2.390 0.425 2.740 0.455 ;
        RECT 1.180 0.255 2.740 0.425 ;
        RECT 2.910 0.425 3.080 0.655 ;
        RECT 3.250 0.595 3.420 1.375 ;
        RECT 3.705 1.205 3.875 1.895 ;
        RECT 4.105 1.445 4.520 1.715 ;
        RECT 3.590 1.035 3.875 1.205 ;
        RECT 3.590 0.425 3.760 1.035 ;
        RECT 2.910 0.255 3.760 0.425 ;
        RECT 3.930 0.085 4.100 0.865 ;
        RECT 4.280 0.415 4.520 1.445 ;
        RECT 4.695 0.595 4.865 2.105 ;
        RECT 5.035 0.890 5.205 2.275 ;
        RECT 8.360 2.105 8.655 2.465 ;
        RECT 5.395 1.615 5.810 2.045 ;
        RECT 6.345 1.935 8.655 2.105 ;
        RECT 5.395 1.445 6.175 1.615 ;
        RECT 5.410 0.995 5.835 1.270 ;
        RECT 5.035 0.825 5.255 0.890 ;
        RECT 5.035 0.720 5.450 0.825 ;
        RECT 5.085 0.655 5.450 0.720 ;
        RECT 4.695 0.485 4.915 0.595 ;
        RECT 4.695 0.265 5.110 0.485 ;
        RECT 5.280 0.320 5.450 0.655 ;
        RECT 5.620 0.630 5.835 0.995 ;
        RECT 6.005 0.425 6.175 1.445 ;
        RECT 6.345 0.595 6.515 1.935 ;
        RECT 8.170 1.875 8.655 1.935 ;
        RECT 7.435 1.495 8.255 1.705 ;
        RECT 8.085 1.325 8.255 1.495 ;
        RECT 7.025 0.945 7.335 1.275 ;
        RECT 8.085 0.995 8.315 1.325 ;
        RECT 7.025 0.730 7.230 0.945 ;
        RECT 8.085 0.905 8.255 0.995 ;
        RECT 7.515 0.750 8.255 0.905 ;
        RECT 7.475 0.735 8.255 0.750 ;
        RECT 6.685 0.425 7.150 0.465 ;
        RECT 6.005 0.255 7.150 0.425 ;
        RECT 7.475 0.295 7.765 0.735 ;
        RECT 8.485 0.585 8.655 1.875 ;
        RECT 7.935 0.085 8.105 0.565 ;
        RECT 8.355 0.255 8.655 0.585 ;
        RECT 0.000 -0.085 8.740 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 3.365 1.445 3.535 1.615 ;
        RECT 4.285 0.765 4.455 0.935 ;
        RECT 5.665 1.445 5.835 1.615 ;
        RECT 4.745 0.425 4.915 0.595 ;
        RECT 5.665 0.765 5.835 0.935 ;
        RECT 7.045 0.765 7.215 0.935 ;
        RECT 7.505 0.425 7.675 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
      LAYER met1 ;
        RECT 3.305 1.600 3.595 1.645 ;
        RECT 5.605 1.600 5.895 1.645 ;
        RECT 3.305 1.460 5.895 1.600 ;
        RECT 3.305 1.415 3.595 1.460 ;
        RECT 5.605 1.415 5.895 1.460 ;
        RECT 4.225 0.920 4.515 0.965 ;
        RECT 5.605 0.920 5.895 0.965 ;
        RECT 6.985 0.920 7.275 0.965 ;
        RECT 4.225 0.780 7.275 0.920 ;
        RECT 4.225 0.735 4.515 0.780 ;
        RECT 5.605 0.735 5.895 0.780 ;
        RECT 6.985 0.735 7.275 0.780 ;
        RECT 4.685 0.580 4.975 0.625 ;
        RECT 7.445 0.580 7.735 0.625 ;
        RECT 4.685 0.440 7.735 0.580 ;
        RECT 4.685 0.395 4.975 0.440 ;
        RECT 7.445 0.395 7.735 0.440 ;
  END
END sky130_fd_sc_hd__xor3_1

#--------EOF---------

MACRO sky130_fd_sc_hd__xor3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 7.965 1.075 8.375 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.661500 ;
    PORT
      LAYER li1 ;
        RECT 7.145 1.445 7.725 1.615 ;
        RECT 7.145 0.995 7.315 1.445 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.381000 ;
    PORT
      LAYER li1 ;
        RECT 2.320 0.995 2.955 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.210 1.005 7.625 1.015 ;
        RECT 0.210 0.115 9.155 1.005 ;
        RECT 0.210 0.105 1.695 0.115 ;
        RECT 4.180 0.105 5.140 0.115 ;
        RECT 7.200 0.105 9.155 0.115 ;
        RECT 0.210 0.085 0.315 0.105 ;
        RECT 0.145 -0.085 0.315 0.085 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.390 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 0.820 2.045 1.070 2.465 ;
        RECT 0.545 1.440 1.070 2.045 ;
        RECT 0.545 0.925 0.860 1.440 ;
        RECT 0.545 0.660 1.050 0.925 ;
        RECT 0.800 0.350 1.050 0.660 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 9.200 2.805 ;
        RECT 0.300 2.215 0.650 2.635 ;
        RECT 1.240 2.215 1.575 2.635 ;
        RECT 1.760 2.235 3.355 2.405 ;
        RECT 3.570 2.235 3.975 2.405 ;
        RECT 4.145 2.235 4.475 2.635 ;
        RECT 4.810 2.275 7.905 2.445 ;
        RECT 8.315 2.275 8.650 2.635 ;
        RECT 1.760 2.045 1.930 2.235 ;
        RECT 3.805 2.065 3.975 2.235 ;
        RECT 4.810 2.065 4.980 2.275 ;
        RECT 1.240 1.875 1.930 2.045 ;
        RECT 2.330 1.895 3.635 2.065 ;
        RECT 3.805 1.895 4.980 2.065 ;
        RECT 1.240 1.325 1.410 1.875 ;
        RECT 1.645 1.535 3.295 1.705 ;
        RECT 1.210 0.995 1.410 1.325 ;
        RECT 1.240 0.865 1.410 0.995 ;
        RECT 1.240 0.695 1.810 0.865 ;
        RECT 0.300 0.085 0.630 0.465 ;
        RECT 1.220 0.085 1.470 0.525 ;
        RECT 1.640 0.425 1.810 0.695 ;
        RECT 1.980 0.595 2.150 1.535 ;
        RECT 3.125 1.325 3.295 1.535 ;
        RECT 3.465 1.695 3.635 1.895 ;
        RECT 3.465 1.525 3.995 1.695 ;
        RECT 3.710 1.375 3.995 1.525 ;
        RECT 3.125 0.995 3.400 1.325 ;
        RECT 2.430 0.655 3.540 0.825 ;
        RECT 2.850 0.425 3.200 0.455 ;
        RECT 1.640 0.255 3.200 0.425 ;
        RECT 3.370 0.425 3.540 0.655 ;
        RECT 3.710 0.595 3.880 1.375 ;
        RECT 4.165 1.205 4.335 1.895 ;
        RECT 4.565 1.445 4.980 1.715 ;
        RECT 4.050 1.035 4.335 1.205 ;
        RECT 4.050 0.425 4.220 1.035 ;
        RECT 3.370 0.255 4.220 0.425 ;
        RECT 4.390 0.085 4.560 0.865 ;
        RECT 4.740 0.415 4.980 1.445 ;
        RECT 5.155 0.595 5.325 2.105 ;
        RECT 5.495 0.890 5.665 2.275 ;
        RECT 8.820 2.105 9.115 2.465 ;
        RECT 5.855 1.615 6.270 2.045 ;
        RECT 6.805 1.935 9.115 2.105 ;
        RECT 5.855 1.445 6.635 1.615 ;
        RECT 5.870 0.995 6.295 1.270 ;
        RECT 5.495 0.825 5.715 0.890 ;
        RECT 5.495 0.720 5.910 0.825 ;
        RECT 5.545 0.655 5.910 0.720 ;
        RECT 5.155 0.485 5.375 0.595 ;
        RECT 5.155 0.265 5.570 0.485 ;
        RECT 5.740 0.320 5.910 0.655 ;
        RECT 6.080 0.630 6.295 0.995 ;
        RECT 6.465 0.425 6.635 1.445 ;
        RECT 6.805 0.595 6.975 1.935 ;
        RECT 8.630 1.875 9.115 1.935 ;
        RECT 7.895 1.495 8.715 1.705 ;
        RECT 8.545 1.325 8.715 1.495 ;
        RECT 7.485 0.945 7.795 1.275 ;
        RECT 8.545 0.995 8.775 1.325 ;
        RECT 7.485 0.730 7.690 0.945 ;
        RECT 8.545 0.905 8.715 0.995 ;
        RECT 7.975 0.750 8.715 0.905 ;
        RECT 7.935 0.735 8.715 0.750 ;
        RECT 7.145 0.425 7.610 0.465 ;
        RECT 6.465 0.255 7.610 0.425 ;
        RECT 7.935 0.295 8.225 0.735 ;
        RECT 8.945 0.585 9.115 1.875 ;
        RECT 8.395 0.085 8.565 0.565 ;
        RECT 8.815 0.255 9.115 0.585 ;
        RECT 0.000 -0.085 9.200 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 3.825 1.445 3.995 1.615 ;
        RECT 4.745 0.765 4.915 0.935 ;
        RECT 6.125 1.445 6.295 1.615 ;
        RECT 5.205 0.425 5.375 0.595 ;
        RECT 6.125 0.765 6.295 0.935 ;
        RECT 7.505 0.765 7.675 0.935 ;
        RECT 7.965 0.425 8.135 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
      LAYER met1 ;
        RECT 3.765 1.600 4.055 1.645 ;
        RECT 6.065 1.600 6.355 1.645 ;
        RECT 3.765 1.460 6.355 1.600 ;
        RECT 3.765 1.415 4.055 1.460 ;
        RECT 6.065 1.415 6.355 1.460 ;
        RECT 4.685 0.920 4.975 0.965 ;
        RECT 6.065 0.920 6.355 0.965 ;
        RECT 7.445 0.920 7.735 0.965 ;
        RECT 4.685 0.780 7.735 0.920 ;
        RECT 4.685 0.735 4.975 0.780 ;
        RECT 6.065 0.735 6.355 0.780 ;
        RECT 7.445 0.735 7.735 0.780 ;
        RECT 5.145 0.580 5.435 0.625 ;
        RECT 7.905 0.580 8.195 0.625 ;
        RECT 5.145 0.440 8.195 0.580 ;
        RECT 5.145 0.395 5.435 0.440 ;
        RECT 7.905 0.395 8.195 0.440 ;
  END
END sky130_fd_sc_hd__xor3_2

#--------EOF---------

MACRO sky130_fd_sc_hd__xor3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hd__xor3_4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.120 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.246000 ;
    PORT
      LAYER li1 ;
        RECT 8.525 1.075 8.935 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.661500 ;
    PORT
      LAYER li1 ;
        RECT 7.705 1.445 8.285 1.615 ;
        RECT 7.705 0.995 7.875 1.445 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.381000 ;
    PORT
      LAYER li1 ;
        RECT 2.880 0.995 3.515 1.325 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.120 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 1.005 8.185 1.015 ;
        RECT 0.005 0.115 9.755 1.005 ;
        RECT 0.005 0.105 2.395 0.115 ;
        RECT 4.780 0.105 5.700 0.115 ;
        RECT 7.760 0.105 9.755 0.115 ;
        RECT 0.235 -0.085 0.405 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.310 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.120 2.960 ;
    END
  END VPWR
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 0.695 2.045 0.865 2.465 ;
        RECT 1.535 2.045 1.705 2.465 ;
        RECT 0.695 1.455 1.705 2.045 ;
        RECT 0.695 1.440 1.420 1.455 ;
        RECT 1.105 0.925 1.420 1.440 ;
        RECT 0.595 0.830 1.535 0.925 ;
        RECT 0.595 0.660 1.605 0.830 ;
        RECT 0.595 0.350 0.765 0.660 ;
        RECT 1.435 0.350 1.605 0.660 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.120 2.805 ;
        RECT 0.275 2.135 0.445 2.635 ;
        RECT 1.035 2.215 1.365 2.635 ;
        RECT 1.875 2.215 2.205 2.635 ;
        RECT 2.375 2.235 3.915 2.405 ;
        RECT 4.130 2.235 4.535 2.405 ;
        RECT 4.705 2.235 5.035 2.635 ;
        RECT 5.370 2.275 8.465 2.445 ;
        RECT 8.915 2.275 9.245 2.635 ;
        RECT 2.375 2.045 2.545 2.235 ;
        RECT 4.365 2.065 4.535 2.235 ;
        RECT 5.370 2.065 5.540 2.275 ;
        RECT 1.875 1.875 2.545 2.045 ;
        RECT 2.890 1.895 4.195 2.065 ;
        RECT 4.365 1.895 5.540 2.065 ;
        RECT 1.875 1.325 2.045 1.875 ;
        RECT 2.370 1.535 3.855 1.705 ;
        RECT 1.820 0.965 2.045 1.325 ;
        RECT 1.875 0.865 2.045 0.965 ;
        RECT 1.875 0.695 2.365 0.865 ;
        RECT 0.175 0.085 0.345 0.545 ;
        RECT 0.935 0.085 1.265 0.465 ;
        RECT 1.855 0.085 2.025 0.525 ;
        RECT 2.195 0.425 2.365 0.695 ;
        RECT 2.540 0.595 2.710 1.535 ;
        RECT 3.685 1.325 3.855 1.535 ;
        RECT 4.025 1.695 4.195 1.895 ;
        RECT 4.025 1.525 4.555 1.695 ;
        RECT 4.270 1.375 4.555 1.525 ;
        RECT 3.685 0.995 4.055 1.325 ;
        RECT 2.990 0.655 4.100 0.825 ;
        RECT 3.410 0.425 3.760 0.455 ;
        RECT 2.195 0.255 3.760 0.425 ;
        RECT 3.930 0.425 4.100 0.655 ;
        RECT 4.270 0.595 4.440 1.375 ;
        RECT 4.725 1.205 4.895 1.895 ;
        RECT 5.125 1.445 5.540 1.715 ;
        RECT 4.610 1.050 4.895 1.205 ;
        RECT 4.610 1.045 4.890 1.050 ;
        RECT 4.610 1.040 4.880 1.045 ;
        RECT 4.610 1.035 4.865 1.040 ;
        RECT 4.610 0.425 4.780 1.035 ;
        RECT 3.930 0.255 4.780 0.425 ;
        RECT 4.950 0.085 5.120 0.885 ;
        RECT 5.300 0.415 5.540 1.445 ;
        RECT 5.715 0.595 5.885 2.105 ;
        RECT 6.075 0.890 6.245 2.275 ;
        RECT 9.415 2.105 9.675 2.465 ;
        RECT 6.415 1.615 6.830 2.045 ;
        RECT 7.365 1.935 9.675 2.105 ;
        RECT 6.415 1.445 7.195 1.615 ;
        RECT 6.430 0.995 6.855 1.270 ;
        RECT 6.075 0.825 6.275 0.890 ;
        RECT 6.075 0.720 6.470 0.825 ;
        RECT 6.105 0.655 6.470 0.720 ;
        RECT 5.715 0.485 5.935 0.595 ;
        RECT 5.715 0.265 6.130 0.485 ;
        RECT 6.300 0.320 6.470 0.655 ;
        RECT 6.640 0.630 6.855 0.995 ;
        RECT 7.025 0.425 7.195 1.445 ;
        RECT 7.365 0.595 7.535 1.935 ;
        RECT 9.190 1.875 9.675 1.935 ;
        RECT 8.455 1.495 9.275 1.705 ;
        RECT 9.105 1.325 9.275 1.495 ;
        RECT 8.045 0.945 8.355 1.275 ;
        RECT 9.105 0.995 9.335 1.325 ;
        RECT 8.045 0.730 8.250 0.945 ;
        RECT 9.105 0.905 9.275 0.995 ;
        RECT 8.535 0.750 9.275 0.905 ;
        RECT 8.495 0.735 9.275 0.750 ;
        RECT 7.705 0.425 8.170 0.465 ;
        RECT 7.025 0.255 8.170 0.425 ;
        RECT 8.495 0.295 8.785 0.735 ;
        RECT 9.505 0.585 9.675 1.875 ;
        RECT 8.995 0.085 9.165 0.565 ;
        RECT 9.415 0.255 9.675 0.585 ;
        RECT 0.000 -0.085 10.120 0.085 ;
      LAYER mcon ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 4.385 1.445 4.555 1.615 ;
        RECT 5.305 0.765 5.475 0.935 ;
        RECT 6.685 1.445 6.855 1.615 ;
        RECT 5.765 0.425 5.935 0.595 ;
        RECT 6.685 0.765 6.855 0.935 ;
        RECT 8.065 0.765 8.235 0.935 ;
        RECT 8.525 0.425 8.695 0.595 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
      LAYER met1 ;
        RECT 4.325 1.600 4.615 1.645 ;
        RECT 6.625 1.600 6.915 1.645 ;
        RECT 4.325 1.460 6.915 1.600 ;
        RECT 4.325 1.415 4.615 1.460 ;
        RECT 6.625 1.415 6.915 1.460 ;
        RECT 5.245 0.920 5.535 0.965 ;
        RECT 6.625 0.920 6.915 0.965 ;
        RECT 8.005 0.920 8.295 0.965 ;
        RECT 5.245 0.780 8.295 0.920 ;
        RECT 5.245 0.735 5.535 0.780 ;
        RECT 6.625 0.735 6.915 0.780 ;
        RECT 8.005 0.735 8.295 0.780 ;
        RECT 5.705 0.580 5.995 0.625 ;
        RECT 8.465 0.580 8.755 0.625 ;
        RECT 5.705 0.440 8.755 0.580 ;
        RECT 5.705 0.395 5.995 0.440 ;
        RECT 8.465 0.395 8.755 0.440 ;
  END
END sky130_fd_sc_hd__xor3_4

#--------EOF---------


END LIBRARY
